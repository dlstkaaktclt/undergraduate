`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dPt5E4AieGCEt/K66u1/rHhPwZDIYuKJwNBuR3AyvXP3DLERa8PZqI33iFD5YJ9K/pk84GsX6gXR
MC76HtZRQg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ipv6ffnwFF7w6Ljnhr7VoRPZgB1xYGVDBO+TeyA+ahu9o3WI4B6MbZL7+nv2IMUuMck+p/96Vm2S
2AlMDXC4nTIaPKSBgF9dXv+35lhtJCWo4bWiW8wYuCs9hpcTZ5QrDse1NwpDrsU1BdGGANPzkO/m
NZcFX3LChIZ7REQB07E=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UZUgdCuw/Ac1ONRQBUfK5aNtN1l1cOReTrgn2gb4ILBz0ZwK5khLM9TWNLMXkoMo7N7PTJ8qzO1k
t50c0i5imhdgTF1vLgLjhrJyhVV36LJbQMbHnsVPNdfrxDUcaUyM4wnvK6amvgGTvU3jGiq3Vw1b
ftPQEstmyIqMvIoyTDwpS5g78tGtVvAxw/I1Du998pj+WRr6NPmYQyZPIzjYyMnEtQCmZd845S+l
jRux0/v8Nl7jeiQFBa5x1XY1pPSUVSaOqNHH5i2VyB4fQGhununoLlUTP8GCP6eExGXfePBOQxsN
5yUsIKgx40ND3sb317vZbUn/6KPB9Jp9AmevmQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
itAx4PFdHKd1pmYBAUAeYLzpD2P3lq3ovIMewnbIZEMg4IhZggNF6oYRG0yDOH3jUWBXfp0UCUlQ
TjLuruS+58ta9malWIYG1Vp2JR7IDWwT+zqneaXOYhFidduDVHGoVSS0s5LW6JITUQB1VxOfbdzG
2Nak8LjI/GUlGwcxphtXykrL89CimAoCE6rE72zVZ0ljifKC+6j9c2d2GMFMUUxIkCion2/IMeT+
LYa6L9Ccs4b2iLDyFdRni+iaXjKg4y7dD7JJ2aKy65TA1KF06xjDS2FxRC20TC1c9JRa9bgaEHWM
oRHZBvkX8S1Wc0DMZS99iNKpcOGPgtcJRLeMTg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hMRQn17JrfkggLuUDBtw0SSucCOYDsiTT49JuhzF7AXT7ldqRnzU79S6QcX2P5xPeSQD1OLrxCMl
P4qRH5kCvfUjpu3u4hQjUZWcXU3Uc8dGpFXYujAE4p5/nCUgMFdnPeqqYENSvOg+CFHRWsucjcRH
dwVo6kCKsn1+vVadQbUqYothaDoMdqKpIfERwVTbk3zbmdnBuq1keVYYsTRE7FewU5+yj0tSQoTG
hXBr3oTfE+RB1x1X5A59k+Lil/UU0AWYuGRJQD6qgv+JatF4ch12k+jUCQWDuKE6qAv2P7aHp5Ai
evj0iRNJXk7I28xo7R+4IIoLSrtcMXVN2rrkdQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
oeVfoBxMjOQlLHahMvbBt9pCmBLpFy87hhFGDJKOlXQpdYbWDCKubxm3l5LJe578FTxJNOLt+DM/
Twrcb4yTwW5J1Ps58huSXu5X2oHCMw5H9jY/GNpPPjViet4YtuG23G+dS3SoW7WoOCiC5XH7F5H+
T8m6V5PyUqGIFLFRr0A=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JygHOAa03zUR1c70sqKmG58tH0oRsKYKnGmP6aNoXz1lyVhXSQACXpOn1c55aV5MmzZUVQBCWZyn
3HUdFXCgloQcywkYOpiV6acnlDrNNZjnJGQkLOmPm4ZmNPxuVGPIZZQtHoT5QUkjbdwDBDPy4jiE
CskQPt97etE7I4zl5d/nG7dX1I4SxKvdHZZChBS/+l85X40Jk3TmO6YAkGszEdNetanqnZZjv209
n8+16TD3e6CyjDT4Oe/Fd9L7vnNhJXfNzkL2tyAsZMCX4E6PjOSMH8NwNuLAasN03HaDJoiPsrvt
3MctCKl3EYFQBnT3ZCKP2+uLu/zRfBsJzwLu8Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 97712)
`protect data_block
RDaXvXadGQd5ChbqAHy6zc3Qhhg7K20iHu7PeVPdpuNV5KcTqlHrLyeqYevQ29iXgwMIVUPrKpPm
RgrmEHw4IyzJf4woBgsM78GQ7SF9EDDnbZ550fihK8PepdH3nt1cxFooT9Om5v6+W7Tz4tUJGsjz
SN06TOLSj4TR/3TGbwVW736xPXmNdFGVLQ0io3vHG5kD8irLvqohpb/t9Kh628QzBgr33vCYblFv
bDcdWvys7rQy+nfEFPCP+s6vMg3YCJMGrme69gHJKrhCc0Oc4SgaVz37iZ/2XX1r6FnUGrJkrEgh
zVWdTKBn6xGDHYSFODgKX2PktMlkV4K9b1nsnE/TyGjGlPlk6beVnilBiJdDNAgxCg2M7R/VIdxj
pO3nbtX/T6fiNmu2QrMpwBTwcAMs6CQvAPTicE0X+xU2FVqzAM+EWkP2fy34vt8adsxNHEIAWf44
+/Qpdggi61pBNaRrs9nF25j+GV7KdUowpA8w04xsXnT7L2zWAL/nDQRemODSV7mcd2aSRCDbfpRJ
8HhgnD84t4GAWK/RT5riLuJQ+PktIEhSekAR4qJ5ZxzlZLWKOehh9GD/mSRaJea/zTc586ajzo9k
e7nZvTfmEzCuuaJWia3ZNScZL5T7VnMKDZxtsp4iAx1Y9xwHAG/VPfDi3LGAkTC/cfYb3WM+gv+A
YHpZ6BsLl7crGs6tRle4xnOL1quuCDli7akrnkEu1qhHMkBFr6d3QWiuG3AswHgRRJ85LE0U5Lf2
EgYFOEGFygVXTMMm5O5C1b5+F/dImLgdMwzb6Zk2GrenTK48cjlPHhaGbZkcQDW2p++B4VpGDd1f
2233t6iOIYc75Wf+buI/eXMTK9n2JaTo8R677ybsyqSoXgXf3nuI47dMCUtEF/ad7tdXhoBbGLds
co4tndhCF3G8zGA4hCNN9/tPnmu0lMy8EOlEBvPTgJtDePM8dJmv/sWyI1GZwQ1EMZVdGRNvQNbq
dUzHXckEkxKd2XDMusLkOzPd9UoEi67DtBX251R987MwcrHEb/PV2IE5RWG0QOCNwTTFdUFAUP4U
de3XI4MayY/65TIET1trMNWikzhIJyc5h4qD+koeZPuLj78CmhQ9BYXVTqo6EzGEgeUHYQXkDcq3
3TvlJR+ilAGc8b8vfGmvFaHrS+nj3G2+zy62kDDakgcR0RM87jczGemAMcJIBDqrqsFK+UdyNlUu
m0JGVnBa1VjeRJCBUcGDhUCWeQuyrO4ZcreTGLM68kWaJV5MGGlcsdcqHrkNDDAoZFIghw6nSEUb
zUL1JZ7EgM4VwXUnlvZjgHcpsg/OXwwKOxTlGCuPz+1BNEPU4YOyCLqfhG77ik/Y2Oz8QM5KKlTV
DuDTLkhsw2g5+4wo5Wnen9UXxnxKucuWtqtGZX/psvhPVuRejfJ+0OMg9cdcQQjEyOKeR0ead9Uu
Q8beTBZsgCxm1gTrC+5kBF+wrMQ4AUliVwAzC4p7zK0WEGfWdjRtroNsWFVmAVWiOUKd1rArVEU1
rzY5Qn8ssNJlR5FfjKwvpVSp3hDEeJc6YSt53TX+zkG0Cb5/JGhKlvhO0X+tLdARMCS2BSYlLzV5
AsSTKD7yqqCg4BxpTzo0KFd5C5lR5wKgQI0HpDOpFNt0uf67pGw9o936+eoHN5VUfzv/aIg9MSnw
RRX82kq04lKjp5bAh0lFGYRBILYpHCP7zbfLVh22FnBHDSxmXzz0y+Tq6XVqrDrTfB1f2Nf0CA92
HAq29tpgJSSuIkV2sB8Sp2IzdqemEgy6ZUCscLj2ud6tYf0Ms+4Ffdk5WyT5UQ614g80Z7Gp1rYb
Pbg5newd9C/LIhiUdapZjxR0U1+aSsbx5IVKj2KITzrkUAubnWRRM7tjITR8EjeBtfWLyhcQ0BW2
GLAfef++U5VDn6wtLzXivnqERLHtUDNqloJCOP1U5eXZGXFAsXFoP0JYWSsnKbTAYv511amAjY9l
EZd4zXh4mRSA5lZeKL89TdxRN03vezHLlSPFe92D/+A7ZPjLJkezp6vi74OjUG3pCzomn6BW+hH7
7Dx8rVJxq5P7IKKJIyPBpiXKKa79/rvG9l5l/MOFNbu3Th+qaqVr/BdNZNe+bSbKgxP7NQeB8NEd
uujoT57w9RUvdIiAUJKZ3y6pjjaNmjvo5hOSEj+GKKySDQNYs6hNd8VycjbqsY+syzF5CdbE0QWA
XYJtYnCG64ggondWeUs7iTTQrkNgLGmSVBSAxXa0ruNzcqGjiUUWom+ZOhwNxdSDXbK4aTA0ipGw
L98a3zZwdejPWHeMGrbKFSTHNOCxPhoaXIBMTkJ7zB/4q4qYAFRPHqkTQXDaCgml+M924BvxDWv1
yXldDR00cjtCWI+QClG7oMOFxJNQHfTdNhSBpoF8/AvdkH66MF9aBbnVUT3YK3aKeHTinPExarLW
VG8ZsJUTpMiWV+XX5Cc1jvHMbq1+3UgDrpv+9NVC8S3j6OiCPee6hbfNTB9fb7n4cZvdGwWLTiak
w0Z0zI6Cj5wEu0Vow5BNm8CRn1qT85H6R0xa6B+Q7MZfqQvk1qTR1P85vhH1afmoiasYjt5zLUOJ
GD3o1hYq2Q4elpB80vCpGInHN19UTg+LpUv71KZC2GT8bdvG4bNYuYGbZFghQrS5hGldRbCRizJh
ZX9/q2Mq2M4PP68clmtuUD9bwZjd1/3qU6WZQkijDdd4kxhPegBcN3xnosGEbCSVNq0vaSDP+r2v
oHvr7HFH+TTyXdCKT4rdOXhzX5d+CjH2QZD5YjvnnBV6wzyKXj+OdzzFITaUUnwBLNwJ9v5Nzup6
vBMO+bsNx35d5aT2VtolBuxWs0c6n5Iq6uV++dEdoq6Eg8RhF9CCmotAKXoRXADYg1PQg0IL8m+q
ED8iN10iSzqC9s4m0WIFyOvDxPGlSqTJoCjTRlCNxZQrwz/AAO1uiD/j0vLJTNCg7aGCKxIj7DuO
keK+sjLPCaPmc9BPaUY0VqxO31rKhEjC9IySuOBUnc3bBo4LDGBNikGa8q9nfjKN5geoxXXPS8Wr
H+RYConh4jEao7pXfyVMtu5si7Q0FT4eKW9pnYU3e/iq7KWHb/ECEYStvFy3oLPIDzwZ+wAoQZL/
eX9ndD50EvsLWBXnx7+rmcgKuSPG+KlLidZ6ZHOSrq39+zIgkxDWN90eyqDebUpKr4JXS8T7jng0
0G4QX88qcVrZOrz5lfRuv21799/J5DK32cEzndfNb8nhXZfcuPy0irOP3FFuR1/w87yajkEspS/Z
QFcAZEuQMcgeJRSUbzBMu8shpPkOEKmV+khbyk6oyLO22TMLChpqtxumJCOvUCxOZZ4ZFMFNuv6f
5g9Xz7M2CsqG9VY5O4zCQuBPQopOa7kDPQksg4MAq2dIxsob5zQzN0zCoL5khKvCyzZNhaSdZeDV
FbCogBa5RDYWrqXv4de9DCueYPoLYujZdw4kTp3XUZ+6ekD8Dfnz4cwzu2+bKavZXskYR+qjtekX
NPpXj1gBGkthC2TmBWy2NyMdo5QKY8qwt/w+j/j+v25MYnQLTB3VVNv/hBIv9sHFG+48QY00nC8d
DeV1hn11Qbqf6tWoCxCMkbVoKO96WyI+MLnK9RqidsxkFoWIPhWJWBNqU1GXUWDRTQ3YCd2lMt1F
Ns7nbhl4yaZtVdJZ+ilJVT5M3BCf0Ycb/II7oq0lgwwHfqBmHLFMNlBNn0oXp3Kivbbvs2u1xOMw
10MmTYPXvbUXz043q4syjIA2elhf/XYZPt8//SDKsbPDSLBQSYwiqfUJ+aBJkwCQ9V4+w8zReAcS
dORfvxZIcLLyPLE0FgXCk6RuUz8z8x614kM3NJk5+NIadOdAiMYpLJQwOba1Lt7LpUqglEd4VlGr
aXKPGf9Abe2vCOyltmhGUaaD5qH/zJ07MEU7aqIPt5rSQLTld5o9EFWmdxW2GfLVksFt6+78r7L7
KG4FKVT8EAG4uNX0Ccjxaia50DAGHdZItYgOnz5ctYj+wQQUExpN4IXKBzmMAx7V+WpON8xfnPk9
aUHY/zNcybxqio3DHGzZ3v16sZeWYPmmOaiVBY8YniIGBx2c616gUkcO6WDjwAM2EZsKMtwoLBE2
cTz1fLmJ3YchRBWdC22NHVneNhm1ZVGPMIxcdd9klg1rcex0ISzopxEatXPX6Q/ZQe37JVje2qSb
KySShwmzW+yNCwRSP/lq+gke3qmcx237QxxCQa2ILPhQi/gmzv0tspN/IMR1RzhbIsBf6rzi0idM
blegQwOHUzmbE+N3Dzf+LLdDtwhbVXqljiBEir6WC6tISal8gWgbyLKIo2of/c8YuLEfktwCanV8
YDEjSAxKANis9BafpV0XCLgwiLQxrK69hkw6eByvQlCZLNFT1yP7bPEy4q10bwfo16PpFAkFrx3z
mhgzpVZ9CjXT4WY/NTNUqSx3jOZv3QAoxSCH4miOMtOdtFl4Qo/uEySZuZ6XSmJOdUeFuznI6OTU
fIvA+QUCJvKHGu0zAwe0x2s2QJr3kKwsUe+gqLzs/As9MQpTHQRG/jn6mMaQtfcmbNyrSfYJ4DSv
cLfZi5eM4yq6rQyz+QlOmVBo9fIejRo28IQvQ47gTq9J7Y8mmwZkJyz7mgk/uATgLERim1niaklJ
qO8sLXeEPKOtpwQYBbjjMcvD2UyP9kUt12YcKbbRz6EUBaK56UF0JAx9xlAMobcM33v2fMSZHdAm
IuIOP2KorMVpAbs/yX2FfuQYOGRaSyYYumwjH5uslFL8ctlqEoUy4GW3zWo/x7apq2WqhuxkGm0t
+U4izM3WhpRLDxjxDPeCU5a7GvUtryY1X8qU4fKgBlURB0UOxGa2cvQmm69Splp1h2pR95cqYvRp
8+nuoxtfzaFj5s+SZI/wFM4brXmOsBFG5V4M+J75gQoflEfbOR77HmM40YT99+6tUj1N8mQAN3rd
a9TPv1MF8AAUrVA+DnQBGHUVfULL7S0oR/N0qymuDxjsbY3in7zCB9HJEb3HuB7i33qxYsBXedLt
Q224Spw2v3hxDW+YxtyJaXKNP6dyKPpRVtlTYpJdss0LL/B52hdB1nWEYO+TfLAar0fJJy5LXeS1
mbIBaF9MIFwYVEfL0/aDYhfqiKPWcNDlhrLL95YaNV+tlKzZ5/htVa9rfUu91PKAGqBea4S4mx8D
EcgQu0BNjBipAYa9AS6c8ouD7g6Vcgcy9bAg/yOFidFCqgu64qjW2ucGUGtEAV+Jktrfj0cqTWtO
GjW17EpHyHTV9wPOLdQ4Ijc6ZnS+UL6JoslAJ2UbDza7ZxtQl1cp30/24AqoaK4Ui3AUgWQtJ5zV
OSAA196l6DcfQEzQKNKiqu6qNbzoI0+j7LV/npRLKiUoxXWP+sMiJUFWzJvuRuwUyGgIsV0iM0A8
er918DisV+0Gme/SmtJNJ9e0LIBzWU/5Rt0jKYodRh7V0ltVh0MYF4/1sGTM90yTDkWBIyD95Qww
+c9IlpLcwBjvLTyQSJq+Goz3F9cAHcqky9JggTDp+I0D5uB54z7zFzQot74sAEqYdN49GrEyM/6j
Kffy7c9wxXxTJjTwOu/FXEUTcM/OO2ugO6G4TddVfyXlyrXivM8H+A+YIAagw0IeZwOJwoq9LNu4
ON7DxpfGjzYuW7Mxlu4nwevlFEI/7EyMrqfFZOHMFlJCNLe5CoqgkmvvRiXuy4Wm0+A7fjA776XO
JjJeR/ysPTNWn/4twlgC32leX1XKj3UhpRRMi9cx6Hzw5xZKoZZjX7Z7CTmxxi1jlV7UCTxCsZwG
ABGkcvtccsE1TNsARd/eOClqgpOW4Oz2VeYRkT4qsfMeprMjcW24m81FeQWGL1lF++oAEFQF78Y7
fWTgW9B2OqbAB3oPBjt+1f7H7kkoWUwgp+lWuVjRQdE7DhcGP677MDh7UNUYfMVEjynfgE1wwOYH
oGy3fmjH7fRUTWTPl6z9shKMy4wKpak+b/uNWq4JPdonimmY3Og/afNveff6dWQSKmy1qzEYg9w7
H/44T+Jw2Zi2JBJoJP09AWI7HrUCxXQgM39BaixdEbFzCLovFbYIy7OrCjjvWhgPQs+jYTFHCmCU
oR37KuHvhmemTF5gP3KF+ligy7vAOwwVsaUoDo5JN/Hay/9p9HHaekKVQjNATcoVmYaZIR4weIFp
TJiTYB1rCqzDcsbqdfMlEWvTuCuSY2DbZ9oDlqyIVwafmW1jHeL+V6URS6PX8V92SszkmFbbXPp5
4fCrGnr4BwA7CrfA/0iACaKIysXfvsYNWgRbZ582H7Pgup3OcwXqIFE0Mc/6r9XBQHg6KvjeCcyf
smssAuI7UioZwFINYb5+Ppah/fadxAm+uLOC2fAnQsRkway4JDRdNNvA7VjVgYnjA/wGMVne4kwo
f9exwxWkeN04r299PqeEQ9feeMZTOwivjWC7ikTNU1kOQ3+Mf7vo0pfGSCOhpnxx2sl7bvs0dKEa
qP/NY8lSgGMnfpK3A/t4SQ5mQigBTerOUYo2bA0lpoZjJS8jk+IfvxSpfKUNhrWRLf3o+MfTFlBo
p1tZY06q3rFFNGZtxjVkfHll7nK9siy6n7sn1jeol9mLk9iT/Cb7TJohsghzGgFeqY3remBzA1ur
Jm41Toqx7/eUhq+QlvNpSvSBj3NzlJjs+7L8VG5fcHC70jktvwmvSk9k2VfGsbJk58vcxYOL8DSq
1O7VOCGuDSEJmIORmrOa34y9NL6YmuzASxm32XBG0+hkuJxhzCjD4ce5T7Mo/Lmbg1bWsYKPqyb2
u6XdkU64fZRD7WpwuUP+BxiVqKbImxvTCJDrdNKfRV4j7X7/dt2OmdA5Zr4dfXYmo7Ro6iCsNHfD
ZS/NgoEjmEDir4VsLW1MQ5AD1WUl5yrkvOMiMq209VBHpctTZ66+A13SNpRkrU1zkxYQB6O9rSXo
pSICAhZl5kgER+8b09CBL2PbomIJHUZhOa2tvZxNW2JRpY8AmNJCmD7MKQmNcyFDYvh4+zzbXgOJ
Vg2ivHxDY3P0nbkO62AJ8yuoRiGEBAt4PNN6tNrds+ZXxWds6VieN7eQ3TXfSHG1i/8c88NxPvjq
9GV27Oknl2waA0VcF/5UCRQDbef6vizo71crirvBaamFdgym/gqWXqeKc/xrng9xZwNFW8SaNPtU
tcfg8llqjy9ISD4BzN04dYLtKUi/hn1gaoqJ0RWTdW+hVY0CVrNv5TPJG3odtXA73CHRLSLKlJm7
ALe+tbMy+RSkGfFo9bsSLMZOTHLay0KR4NJ4QpdjoXhbqFC4BDR5EUcS9cnsmoY9m36bYbbMl/SM
mf/s51dwJg2UK6aX/+8MUM6jhFm6TdALd+KIj+7TsPV1px4cwsKOSqKd0Scr1xzCyo07sOQ/cMHX
KYZMgyfZTs5tHXzNrzkF/lrsZl7zwNeMbfa4EHBZGUYxe6YYEULnH1keFe5hv+xUhaPKQqvPsDsv
rv9aTwCB05s5Kzu4EgWAYWd8hxCdN/JU1PxVb0XE99SEL4u2BEGXhMqu+lJuHj8b24fG3B7uhIEu
1IP5cLgT7754FSfAt7L+usS9YvSXsJyaI/l5lMhy0WYZvC7dVAb+BAu5NWVCh9N9qq5ruevZkyfk
L/P6NBnRPVDMO1a0/NScd9zUL+OQSBfapQtx9NT7hedEG6G3VHCtnI941zlrWqNPPX/o8NoUVESk
G1c5QdviI/rIF7LKlLb+WslMfAO7opB7s5X6HwU+VbKuTi+0vOP6pbzmPyXlKgQhDzNjbXvb+BLF
oZbtJ/5CVL1Cv6TmJMJNqMZdWyqCxpKQFH+1Cum43783H43AVFTk/PCZ5rPPQWsqNc/iImrpY6zU
TECsbw33elUSnytUo99u3b65+BNmq7mbJ8xHMqL8jA105dKOTNpPi9WddGtxmmDcyIef2zBPTGdx
AKa6WRuAe2QxkgYrymuXubpz+TFQQoc8a09NWfZP9FKaqXShWMhM9H3h2RyzOV7Op0gi1jMyblrp
vH2C8DyZ+P/x8fn0Ek2n+6eNh5PnlMw3TJdcMMyjArs0vFofgmDFvxABrMafloC3/33/8BfjyjPQ
8yMaIBt0BYH097QAYpSCmHifzoS1l0q4WbyPcunp3zvITeQRTnE7wtXdcHAMddB04NvgnafJ75Yo
hSVhi9QJl/aVS0gSEqMzi/BcKEoRJVRiP1MSegb9ojkyeh8+DDEid+poe1RNTWmJmsiv1xtnh93p
M29hhiS5yqCwWANeM0MvkPLDlE6qu/2uL9A1gRctiArd8OeKL5gwEHUYRwqqrQf308zlZW0XvW4x
AfXqlun1wjC2KPTTIHiMHUYcfCIg0enWxGH/bhaVquVAco07NAWVGHggrlWuvW9UlLLdYGFxWDap
41ughVT6NCGyvoK9POPmPmbTW4W8WgHOB3EY1DDZE1XbiJESz4sPybCYUyM/p/iS24NRjLbs9AYD
yDfRQvMm/lH4BxKhHCMohmZyZfTpEGHdr5qh6ueIYdCONGW/FfZCmCrD7QZDilfTFYrW3h/rtEth
GQZoDJj/404W8KDtbc75uQipzQJtMSM1+3+aADt4og9j/zqtOUrx98AuyGPfAG/FznAsQOvQjGm/
zbpKbNiWXoGXW1XdmkSjkQMMWhFQOJ99rQRXjvHIGK8Gb22H92MUrTpCGiA5nDTjcoqJldco3gWz
3BIQ53Inu8LhVu1vne8hlmFvOFQrP4dtew0dt8nbYXW2EvtZnkwCvggN6i8kJLtAS85d0s9FSOhh
4hxeblqMM7mofA8l5eXdIuqdt9jrqE2ypROaJOMJJnPaPKhDgAA/tmfxnBmaFJiZPfyfQRMK/4Ko
iBrAjtbuCcw2AFQR2ng2Bozo73UvA1GLnFAV5//tvnwJWvgVcE1pJFAZGuu00sZUgXLLITf++6Ed
DH1EAcIunsn/cPgSCjJc1fljs80OjxYqxnDa6KZguXmp7oRcpMvkzfN3dkLsvoDop90QNM2bv68/
sWSQJOCc2fqvIzdQhLdmshsDNegW+WIP79a5TzIjmtiW3cypMOl+a3WsJXcwyrqYsTSIeAqA5RQW
vAjqxoPWkL23aE87wbO12aU/TYPO8Z7+ZsPaYldK40XDjqWwHltHbTgdd/l5ivvrdmlTnlg1yaPU
JXEo1Ry+Kbv7IpIIMKP5tOx+ZebW7hMSvRLFcLt7bOzXHX/dg+h63wzi7dtUBDA4VKrRRbRH49SY
cVv7OCW8hbJ+rpEEtaCdstvhokkHD56opwXTgSnEZ2gefk1iIBZAcn2f6I3ogz5FyIqSHAysVLWD
RqK2GpzU99JzXO9OZtEPrfzPYkLx6BDS8jfxcPREkaKk9sjagI+23ru1D0UPVU7sRBEuheaifvXh
n4ob78Sh+soaeeGD7vr0qcHDBhjCgMfUw5CIQ9aF82YWBVlJZoHKjEu7PlFvlwK2kKovPABsn9eo
rVvNlfDskqGWhAQLw+aSrwa+yabcCCeMis9LEX2crTHjq12/vRI9ZUHiuPfK4AVJoHQo73AejGQb
eeUMDfxhgDbO1oRXI8PMa96oFza7NCmUiO2vj/pszfYCLzkIC4lvrpYaz2QWv4Bdz/Gt4/qYV77J
sEBnKkIfDZnGfEJLWpWH48HwZkBfkF2njfR74OUIPE4XpYo31W18k8/sLjhpCsl4HtzbXZA0K526
UmQ4uewVzedWNpVNdzHTpD+PGMSq7T2QdL+bKJWNWYzhWDfSj73LgL34YEUh+j2tH9q1lmQ2vesP
LeFbEoWwowSblw5Se5hDgepfW7VwTrYisvWQkR7+PWOhNP5rgFwdAFxlQLQkVGrlMgooCuFzicGz
xRYA1JvH2V0f/Ayb3N7agw/GposOxDrRDaFS0lVqCHGvM32RbTVYstna1hObPHaCzkeLmW+E+Tk5
WQpPDXxV+Y8s9N8t1wsR5O8TZ9VlCR6u83Y8/Y4D/rJjrduDdDPCK+Wx0UcSkF2KKyS2Yxpio2US
XYACGkYg7SWa2bqtJ7Tmzne+GztHz4cuVulxrlFcP6hsSE0ZWPYEoatj//n+HpgHIpWr7ZnY/H8D
jz7uHPZ24U/lMYQdzjE5CcjhD0DVd/rqD3hN9uFGvWFEeinWi08xzdPn9OwEbxv46kHxV8vWngJT
ovS3s9uMQng3mL3CdeHRz8mdgdDMmXNfOuvv6ilS3Da8pjBwGCtLMUUK/dIz4R/oDQzfHwBcBpwG
34SutiPzBs9Nhe2TKI9dZ3iuluWZ4tOxeQIfK9jStRWOhgXnrvILkx78edOC8w/cG8UuGtO1Gzj5
dIXl0+erqPOoHh+PsZTRJL/Tcl2K39AFdg47Zoztyvvic8A6PmhzUI9SNckwxgdtPHLlraPCXibd
Vr27o07I4s9/yyZ5KhnBZ3SQVjXmaNxuGEKc9x6gIgyVkVr6yLzCb4BbZ9HPpsydmfvfwJd55p7w
92CdXKE/j6JZ3vH/JL+xZ+Y/r0Mo/fIhtaUs7g7R+gHW5TfB8GdhDYy6XgMN3xV6YjsLtU+2q0Aq
Y/GIvVOyLaCnmYY82pilIYn8NqgcFiHcEIYuW2/aK7/7Nyw9YoeAufS3HLDOO5mIQa2Mg7LvF7nk
De9uenLEz0tr4wZimkKKdjcsHZXRRu2x4neFjse3w3gMkgZ03LqT1Cx7roAcnDAi09ix/2YA6SeK
Dr5Sa6tqHSiL8ai6M7nROhjm89FWSTM0D6hXMwxF4GApeEJC0sBt/geRXtRwuetVX4Akxb48yhfU
U75urY8rkHHANDTDF2D6/kTFrN+0x0C6Dp2rObqcgwXZMjNN2J31CA/bZTwJ9+SEf6NukG6v2KkR
quyeDDOzeCWl0eNlXbwp0UBc0Hz24hG2rgb4/TllRAv8wRXmLR/63QWPi+CC8rJkdKoXrZNWIblQ
/cDFr7Cf2EuQmmYvAfWcPYSYmmvI21XOakkIHGK5aS6gkExRO2ClraFruRG3jgNumAHmXIkAAy9L
TYD7OnCcalCEjs4SlyJF4QUsgvROZeN0Z6cC75okQhjEkY+g+3y6+PvoQyAm7GXcO2GBii6U9uHW
2/9tQ+D297ovLyMKx6SKgOEsh/hgZ0qXnCUIcb31Qx8BwVh7MdlJ8KLjS4JUz4d10aSXzOEtEL1n
LYyhSu46nvGCMXMFbF6ilO9y4nbHFov2GGSJIe4eh6ObuDD+7aMqFnSzowVQIobLvutNpXqK1iTx
2D6aaTlD1Xj7+qVBMUTVNswivjOQy62kG7jAoWbjFpMa1FoT9PY8/5RKpITxIrUSAMp8Y6ZEY/qn
hpm09kFHc9nWwcdEmakIzxYpf7GjMRqkFEhpHPTzRcZOFM/f3BIyDdFQquc31lmvvVVh7RNoK0Um
4STSrXutyP0HrkHK+TKYtJESDk5I3BaPKcVWJmI/KYbCoN5Jj16BvZ77Xg8IbplymUSBs91G43gY
Pc+qfN2Q6gl0InnxaXUFNXcJi506rk+aBn0GXpTtxeLYhor6Cv0fM7XlJ+/nd9twlibvUrPHcDT8
rgCKzp3I7RFFBpFcB6D9nRsCp/qXlId4E2wKS7wR26DRtRulnWIJaGfLb+B+/vngQ3XTv8TvR2vu
MngBQo473AM4OHVZqXD8ykA9Hk480gm7/L7hcFINvx2ZYEv4evw8a04OWIT2FtJQhVTkbDC1DuXt
aoRPB6Pa8+NJzueMvIY38cj6q0TImw/PuD/zjr+2Eym7MLWX0x1QWp42H8taACzTYqpsqlyn1M0J
SPzkQXjCBclHUJOCaHHMK67xvd718Ix6ELxDeS6z6bS4HihEfcqUIAdVTEmf5BcoS3lWRyBByTtt
uvYcDjJJFy6Q4yIvV+qNH4qjK2HWh5CGj5cgbOHT2RXeeiAVa02MZ48w2p0L/xnlJQNLpCPRC+CF
CxiSEIhIfxU4u4hFey1E2oqxtc7Umk5QiEBXTlcIAJEmbDxWuSHjVcTYQOrw1OCC49RQkOq1bWBo
YObAMx+E8Ao8LxShqikrntpV7qHDp6CG4By1inVVxpp2QXonNvsw6hfFD5+NhTRHPGROfnkXOk7o
OFFAFOvWk3ePLWoWPk/O6iSlii6AkcnWMFwGf1v/QceuIBjYJD/xVgdvv3GRBMIDAa10jvWXyrD0
5dd7TPTxwzmYk4VFhJ67saN70lapFMgxxHoSqaAOwUg3FpG+2nU9AKB9NGMx8GwKjeC5YKOPs/7G
m6Tw1z+ORI3DS5muN695zDgAjL5gUxmM7TNf9e98F+nfnD/z4G57Jv4O388kNKWcqaZGqAMzae98
NElfgyWCeLQiiKR6uFRx7/Sz7K+lmfEouXt886hZYn4Vd4fJXe3I5cGawnECiZghQ2JVHcT3zYTN
zlKlSzuNsl1gfkkqB7uwWcyCT7af9+jzpuE1M4d+ZenAoyUSebe3h7f1gnBOcLZfhm2VRkBdkw4a
CZpurPBNees3ndctx34/Ijfy2rT6sEc2rNNqHuLdOGsA1qQoiS5MH4nvZNu/NfVFIXf8DSLgGZ2g
j7UtrO64TJz78WtS7/JnJldPPuriMQX84Ae7bx5ll5dPL+bPobgvggkN73m6yK0vm93axacr0U3z
kKPVuk578/HMtSkrtEifzm1VD34eo86qpbl20bUHM+9BPf2efhzC7JAqt2m2OiLbdH7qkwAKvocY
c4peWkWgWV7pFZPiN3yk+YWYGJjZG1Vf9jAg+a3fZwUWhD/7aBPOnDaAjOahnCKJi+SCSKyCr7+D
WeS/akeu/40am3TCtNoVQ7l0vD7BEVPOLvw4HqTx1ga1fnlkVHWT/cxORak6qzptIyjr0pnfhwSu
ChIKCY3+8l1gY2mjNVwaqASexAVtIkWNU0x2yrSKg39euQaozUhNmjdSeRwL6F8kozLUFKmRcoj6
lDaVBo+t00EXXSZtHOi8OQlz1E13gaGxu4utTeBjR6qre1pQxmVd92aAkluSC13UNu9IqaD+vkU5
cMdVO3YUgNl8ggWO8iH9upMSXY0YoMVVjZ7qLcrn/yyWw+TdhEf30+6cxi/OiO1gmFMpQeMMlA4B
tmspMEZem2wkdbygzmIrhkJBZQ4yvsdFG1E8K3hMSjUS4QfVWrzCP0u1ZNgXiQyRh0bS5eTsUTpJ
5rCc4fK+b6GpV0otdHe+e7vcrYIz0y2MVoKudGdjF8y3eHwlp7901JGKgdq2ixQ70r/Ai/Bc4Gvw
zEIPV26Rp5v7y05yg/OG97dwu72sEGXrpbD6LOSQcfuQ6djcXhzD+mQ4zlZgRvxdg+UL+QAuQU5W
w2ntRU/A63L6GBBi64vFvu9oa/vewM8xANaTHgfgQoBiWHZrXPg84Da+1qQhmfoG+fxM3wQtBEUF
mXg6gP+DN1NPXY9sw5vmx1fF/KB5+3O/eeEC6sj2sz5yzVzpY4MUCNoAbNvnkdGPoyR93xZh2u1S
/Vzts8dYU8OxIzbkgXl9bEJ8xJB6P95malRcFp3tIoSQl8TI1ym7lbeGoeAzn5rSRonjQXunLSHQ
ns7uAI/zv10GXu6uPzlt70iQ4WOt6vQ1bSpPFGPmY3mdR5ny8RuPLGJwA7Lv7kNldxDA84nWZxG/
MKIp2PHwJj+wA8/O/ie/W6d9a5MIeeaBTq8OCkpUxwCnEB0pPJLkJhyt+6dti/Upxk4bpndByN3G
8lCqcpveYP3pafccEcrKt/FqZ5ODyiLxs5aUkia7U6CI8qQLI01w7+L4KlVYl4/kGEflKVpJ5VJW
zjZe6gRKjss/EkMLSBMJQKfSCjoo3prwFoZOAPlrYZWV/YL9Do0FkBEaGHB/TqxHbw7qTJ2u8yYG
xxtz2fbq7BeZZA/HR1rng5SDRP/OGEIbQyG77OC1aigC1IxSJbOlUlXk81I2Pj9hJ23510LMXEjQ
mLa+o7p+DNQRe4J2Jh35qYahkCEjDAYC75+Rl6qplOBQwWFpuwp0BCcm3IHHErv3ZDT+COy2kmzZ
SnkkAhsgx6eq/xKFozRn8pN07EIi6/esEfDIS3/ptcdnMLUZGsc1PWZpC7HXCDgOSaWkGey3qGYL
nhV1vQdnhP82KXiCCAeiDP18xDGybK00ya3JTQfpQze2WaizI8shas4HfoAiCNBeyUb1K3Cbxft5
WfTrSaIYsnYYaPonNY2ULyqWrEgoMCnSK2vzAFuXVCeSBPAJOYY2ALTJem2gX3GtEJUdQDLUqtol
yXHwdWhDQThLRGATum72ZvU3XyBKQrFOLjRFSBhDfhDqABhpPea2itajTWj6eGEIMKVuUGMdgyOb
tONLJy/dkaboH4gzPe8h5DfKYbwrZ3BBKpw+Dw2dVvKl0M+jvVCuQjJb8yzLJ9xQVcg+Gql1abTf
9jWfrE2oFZV6emfgBGmX0lrp4xXDMhq0Xt43+LcikpPPp5M4yO91HD4WYywcMO0e2ISrIS0zbPZK
nmlxzet7idSBeoDc06ZjnGFZwQYU1crPfwk3bX7KdIIM5vOoxKNU46M2kUTIyvRvJanupYLDQjC6
5J5Q8AYA0LTCvis1GUYMl6IGTK5d8zCdzMvOkC44oa/gsvfx8uU28+Gj49K+/ljL2WCrHmE11r3m
9M+icfq6KRddQYAgrDWcYybsHxOmITLCcl2JriglWdnEQUZBET2M1Edgduj2KsVcxy1Ao7Bko6HD
KZ56sctqC3LtgwC7fJVBpfr5yXVMjspSq8uTvrM84cn3YkQ6CtiCK7Izb9/GhBWWerROi2ch/AR0
G0QnyLV+CtiGQ7nYvCUlYl4dN0/lWZZmijTKLKsN+0lgwtVinJbaT18UiSaDWA881vODcd6u8B5B
oI1LeFMaiWizXfC8M7hj5iLtGwfl3eWY0JAEKZsYJkI9jwmKHYJNZCTlNbbE0dUP0m/CBfgWX6w3
71V6IVDFMt1k/ysgUL2KmtB4AHmr/qgXen840M848gkJVaW6FcNXyCbCYtl/1uA7kHHLQnvMkmrd
stFWCkfipscOqiTEettBsZ6LiieVq2boVUiBcFcKszzoieNeX7CfZZatvI0nz6TNyN6O/3XQHAld
uU6Orm1ZzguUg25cL7xvZZhBi6T7wcpLp1nx7iVIZRba0ouQw7cY+lCxf8PCwdABT2YcCpCIGSLk
QOycQOFFr2kl0Fk4aumItuBB86Ujo71f0FxLTljl17RW7y7d+cptUq4FkGfYFHylEYFCEpVAE55s
9vCrD0U0LlSylYK4n5dYpIqRvG1Q/vJo2fpgVSKd2rOuqUB13wDSjMBurvR0ehz7pknENgAq41/m
N1LTlebYJbbk5pNsJ56o5baRC5GRQ0TymUB9Nxh/nE/IMM6Ncl+aZ/wmAN2lKIsGvhnAgtF90Tl1
olE4tabbpR28/eR2iiUQ6wdwzqw97OKrwGmQV8BbH8zhlUOHJ6rg0XLtfekd8sR9VNOKYam3Ikq2
xPulZcw7UkRgMTS3tad+975/J951AS/Nrea0nu0qA2S4jJ9zPbxg6tsABBF+Eo+6kOauiulnuccZ
WtKNmrrXVNtr+l5pd2Sdkzonu7eVY5zIBaZ9EEVYKLRRHFqRxs/WXwzM5ZqpbOUF/2ANu8b1vSiY
ptX11iTXgK1C+7TumvqcnasM6G77JNECySVDKicENTzM3fYW0oQbRqSygK3k643YoIcJVlLqT/cn
YAhLGxXDw8rNenM0CN/M2Rq9gEVqbHeV8FuHAjq25BuAXQEc5vsXDHwbOviRhyint8fqFhLehmsr
NWXe5m8i0ihu8znqSSKWlf4enFVXnN+ra8SPt3LbyLN88bHkUIF8rV9B3175CXI4v7qx8Su8xxzZ
Sqbnb4eCDRUr5EYV5Qx/wkaS0lxEkiylxBfOxee9E5wNPmgOaKja9HjaMzzCj91T0csvvkopsbKD
oQhPv+d5uJWuA0HfJ2Ky1Ywi1t9QOEH5dQ4nItgd2dhjbCS4ivFNBbZl1nePXTN7Lt0K7bknxLF+
/Mfp1L9D/EFtrWkudjgEp3hWLLKtyYX7CCQ7cyfr2zXv/Q0PHmz65VcBRq0D76e7TDkWmuSnB/n1
MYxW30DM65ZilD8p+09XAH7heguwHbzd684Pbq7ljqEGP+ZOVGWXyo+WDGpPB8z+0SKA9axJ/WbR
eAdMKPMDld82s7I82cQadlJY9O3tRUo5MzTQgv3NxQUNO0WqpBSkhS1o4F1rizEcDMemNH7pIqir
5mTVu3xA/FvELPsXTYGEckpD8RABp9iITSqWga7bThbPob44hRJkCpH32/GERLPT4+0JlIT02K30
KBglIBpiA+0HS0HVm4ngK2uk7LxnCjC9u6VG5FJug9qh/NP+PgT4MvTGe20VYc2cjtIJF4R1hV5A
1JSXG0FExCl6mMD1cxqL5aKwPuNmoug2KeQ0cr8o0As1ALuEgmy0xKpHHe5vSi4jhJh8sThi961Z
0jdphaPzmi3yT96foys6D0TtjVylsyIRyYGBO1cUYjId+K8jGLxr/wjAS7nSlG0uaobh55xMeCyL
s8VYa+fPMaLMvMoVi2XUCYqhryjFe75tQTntlOBTMpFd92s4q7p7QfdA2mmBw6rAKwvor0666A0I
kVMyqMBHcbnsrSQZRJqFNSnW0XD0yDCKaoZbicatoTHUfc6Es1vz+hTmooTfqW4Ldjr1IWu4L32g
fFys9b2j8V2Rfxyg8r247lUAl8AgB8lDSXXPIOg9tVJgqTywybpn7/6Z62lx8ZC+fjvPdhPsfysA
8xzj6aMhEb1QWEqjzLgxBB19ijecJZIve4E2Imodm/5PRZHy2COFLL6yXpsFqVw/1v/xacYmQr4O
czhRv6NrF/CQA/OGIAX0C+bJKWtKhF3xy6E4W8rntVTIpD05h/fBMNSM9egNPvKHbPP/vl+caJle
vYr4zPWzgdtOXlbJsuqCa7pkcmlFhbkOVlB20AlNss7xw7AdS6mWUkkmiqoazFiEGsDVNNqy2+J1
kFaox1uCekwkg/hqdMtxM6JuxrlnFb/BtBYk4Ag8W3JtcVzbgVuvDG5ghEQdMnfeU9PNN4qgRktg
xMDMe3EprMV4vJ74hHAIO6/TdZcdgBklr2lPBBg7gfTZkKAr2PKzG1W49qUVGzly5hP41KvgUEJU
ci+dyrUfgKBFYaUfHA8as4gJIA8eVpId0soXJINO4xDuCKP7cg0ao+xFxbn5N8BLOI8V60/x2UCr
O8HkAsQH+oDtbS9PbTOZ5sZmX1BaFISiWNJr0ZrB0sJywqdloGwsg0xrUNn8gV75zo6clPF5zoDy
khF36dVdl25QDvoC0wCmXju0qVJl1bonidIP4GySx0ldXsn1fP01zMScE7d4PUifpRd5AIbyenWf
9p6+u3u8289TjfWnFxtqmGcn9vGBZ7k3SX1+trQiXX/ypiCK0unM2s0gNpaZVIhBDtVDoYgN27ev
BFnRX7LRpdfBs/l7Xbhk1NVUxrDRAy7MZZuSo/lcTwjn63WOtWgsm8gOAsK5BRRp8bqBXaUDysO9
LbpqYe9lp3ieVwVDn/vFe6XxZuHvO2P02VTzfb0iT2QRFQAxYk8hs6TBa8DRdWE6ExbrmNQGxjmA
87z+4LqFoGA1ZV043WXedag6firANOUMZOax0oZRF0REEQ1lzrgbXXRdE6pIL3mDSBhFE+dhdRf5
fHNqF+LwPPyx9RvHMjDDUvXMcsi2aKVTOkcwWNqDClPikr4y5W2f8uVDG0F+GMM2yz+p4rQKM/w2
XKE6BveOSNShm+Nh3ZNj6Wd1W2vDXG1ikHHU79COA+N5CTquuUja4XQoFowZoyhsL0o5oDuTdQ5R
ZQ1xr2zJZdCfESdRlXWaZksihdHkLWX9VWIjSip2gvNB+A06z5yyCwmtUBFH0CXmIwTEmGf5ZPVw
eO6/8+UyPvSekHUN2i5287xOmXHVzC5ebjfIGkbQokS3JOH5pUZ2MWIqnroWUhvulf33pYnALjde
EraReI2+boKT2h9cFErcsjtMblI3HfHS/2tFVBofu4M/Tt0ordxi658nN2+Q+vCkKOpfNsJ5PzUG
EGKNJxebWUmey06DG2MxhHiiRR4ehD+udPc1L55t8W4hOcek2+M18E0l/HVFqk75MZ18XW8yT/Wf
Fduwd0nC78g4hkU9TKJ+BYlotLBvNbMRlwssZuS9LNwarM0DLArnEQ3+KG2DBJa8vkplWflKxZ4r
94UgEnSQy7ZXBCVr4ZNcJgxTBZq4uria1zm2jEpqEPepZ7bUx2OBXk48UvOGtLG8jtqDRO2bWpN8
EIxgQfCIJVXicHM13TF+9mrRS7rg+wFzGj/O4xRJxdIyn/zpSTEHVZy+Ir5wRvxaewVsPK5u74G/
W1FCCc+TgQJZmm+cvu96HflaPBAA7HVGwPycWLwEmprbdqh1tDrHUEryrRTuiACZIxt1Z4i5DtA+
v/F9jCmwr9Z3karK2XVQWX+Ay+IwfUi0tP6qRuyicWlUd8gwyxZ4Thq2zb/3vwIyNN9TXx9k24Iv
XxELqCv23CCwAPT5/U0FgL305E/mapgMEQZheZj/BllUL99ay8V8iiDLRHuMRb/t1gM1de4KAaTe
ovzt/QJn4KsCX84vgCCfVq5qdSYZ/VTmrQe6HXytXeaWxaOMh7iYpsgiNQuglZDc6Q1jBFRbtnQ2
aYCYFZaZuqWX1Rro4HWrbjc90zUc7v2YzQB41a/6lE93aIhPticAYjqK3vWUGr6WBrgSCiJDHe5i
7UB/RYV4PyhPGeD130YMMTRo8znFNDWu8O/I3VksBeQ51UqCCWYg0t5L2rAheYWxGCYnD6V00kjJ
QPk+ZZ7lzXb9q8sH98/YC+o6H9XG/6O5cp0/m/wMO153no3G15FX1Jwkrynh5vI6hfu8rwPyFvKx
ICkXQBlSfp5+7Ykqr5xtpyQBMEZlHo6cwYayez24uN1ELvZDLKp/IHK0Si9ie9/MROaoEnA0wzXw
+YprRCiFYLLQpeYhRp/aR/Us8GruJ8pvCqI75kcKFjdoqHdZ4NzsfzPE7+sKgiBFGV/kmr4x60KP
O3U/nIBOU/4weFwLRi0AlFamkshguvdePNW02EKK3UmtbRO47rO3lSNnRblH1sjHy7krcKPSnug0
UjyQ4pDaDOoJxCnYHK8IZ5tbKwF2ykyw4jQ4A/wGnTKvy3qczeEYF2DkZ9QUMA213Auv5Ve/HiBJ
Oi+5IV+ia+SR98CdfxyDWAIp24z22PBmBTzFPJy2O+bcITOPwG+NLluNupxnKxivaRZ53MK7PpCi
dCTgsBGrGhRg0JzZGuFJsY2D/Ix47a8Zuxh9SykeJ2X5moEhvE6xu9Ra3HFUL177CsnWfwkcCOM6
yjRptDerRHRXUYOp8hWpFVQLAo7D+/sgKo9kX1wVCMUbO0Dul2fxZU9WQCeJPhSd2QWy7jdrDXW4
vb1L5SSnXNBRDgZPSbFmtnjqdVEWjT2wMw6q6QkULIwa8vH0srb6vsGyQStjRQ17GOLpUkYVwlxY
NTN6KPJBVLJVx7z8acB+t5Lxu/LTGMtv+pCAt2iYwfBqDzrqRfIplsjlQXqOtFK7QulUYlTvoHks
fCC2XGwajTacDhu3/ZusGDXqNeZtN0YaYQKa/NI6UUtil4HMq3zeePZvkBAotyob5eH5/n+KoEdP
K8j/L/U9vbOAucvB08/GEN436OqEemqXsumN2YKESZEAvw5hYv8nlco3/bIOoSIWes8FUcTLhB0x
QKkXLNDqmwBxHne0y57ry+d0KdiMb+q/+mVnmKxPl0TIDogarL+0i7zhQmtc+VtzV7whNrM9x6Ch
mBoXy0qJuQT9pP0NZIwaj9m642wMmJrGPuq7ltnVshccJkQePO/a3rzBQz1pm7YlmlrzjomibH6h
l76KbpYbIUEdtFyJZMO2aaROxD3zGWZ2Pxdi9aIfBEir1C2hx6I0mbz4V99uCUJ7jE05RkzBCaU2
kskv6Gqe9x2vkr05XPtz7KXII4dd/D40uZ2JfDL7XnDs/+72mve0bxkZzu9Un7ASOHqH6xbgCLUq
ugKg7cvPhgjxhGV8ZgHVB0qdse4RvpURbK9sbHhD7b9iaLQlLMNkgoMEzvZghBh9CgzZyj3V2JnE
309T++3SiWXO5wZw/0NAzcb4f8qVQIbQ4RGK8DMGT9tj5RUb0Rr40fPZ9IZc4qIDB5UhAbb6eAf1
c1HLI+dqBfb5D2XvHxgBgvMWCUn3Sh7hVh9HRufhPsZwQ6aPOtsf4QhI8IOGJ7wozrXo03TGTaav
7/Jm0DvhGMIWH7/aefFCinOtxruwoqTOHWihx1eboCyW2sA7GT1dPxRaUAjOz/HMsu3ty65uDjWB
/jEtshceo5r+gX85y4W910sJFX3fH42mlleB9G1j9hdzfhOE7dHtWjGhH6ZXYfDItUuSXMG8PGAO
NqgFgG09/m4WrtM9ZK4xtN8c3EhT03gGhY8ALIaSxxywrk3fGxp1EWNSI4OCGc9VZhKDlOT62Ktu
osMdqsLHfc8M/m2ja2aIfhENlgv3Upzj/LRyrVG4nFmLgg4MH0hgnxo3mu4LAwXXOH3wRvMdv9nd
UU6taCH3vjH6Dg1w81fxSaspjjIw6ZSbhMYyHw1zV4i+q8XJbuv/p73Y6ubRzy2E9Psdlb0YMIiZ
b+XTODqpQHoIO55gcUEjZjXniKH+XZc+0w1JX77VBjuxPCYR59adBucdNPRKeTKUTtRljdZuC4CK
Y/+0iBvn0+nVMMB+mxmK/sGGZcWyN4vEGYN3Wzh6SIzEK/Jr6qMl3/5tKlfD03AMD9ki25qEsMib
IY8Javi6XaAqKSTXFd/VuWYvwA3dSz2NQfrJZFsQnUnB+0MLGlTU86kde1KeS6KY4IYIjteIXBR3
xubpXAnEmkRU7LjC53yYJlvgu35igr3WxQXv8nNsU+mvHSIKlPTosBbbcUy8GSjybzRjH3POqCjM
kV4Z2KfFgtn41pUutgIGqsXmu8ILtmmc+aIV0sHYpHzgVAWvIx6pj/KpPrUOySm0+LkZa6gkggV7
Sgq+kL1iY/vQTv5UELkOx/lrevw2rtBAuPeF1dQsEZbncJXr58z7tnpOUJNSyAlpDm7sItg3EDTG
Olrg+Q4IwfJ1kuSf3TcL/SXjvPIDdSVYioAqajJsFc+3jvgfIWlVsaeF8XZMH7WJb96sRIwR9gLY
I1bgyT38aFQj7vqOW08ydF05k0K3TNpVsQIlS70X3XzuFGgLVFCSTT1XrnmIC4csO8x1Zppel2J1
T8OaBWkKjki//+OA8zvPNriVKWMiGAZ9HjGAXVsTBHyDuIp54N8Dnmvu9eKNiq1s4lwek28MfdAz
ldxnZrHNDDMX54f3uzYYKcKi8AgTv2lqmFrvlfo2p8KWuprrA50AgtgCilSIKSXygNOmDWjbIjOL
cWh5zOgr6cQdGxS+tv1/QZknMsoBbLMDOwNAGLMMUksELL8WnvEgFUvI83h03pX1rGjOBf/ZvicW
qDAA9sUAJ0osJTHp+KpNpAcyeZb5UGtwhyH9PveDNAhfQx/F1B341s8ffYkQvKQeeTQ5Syk8plHL
eJuPTLwHDwSQr7s5o1LthG4qCCTjDSUqhzv1jP8LF/Bc6Qy/G2aArC9v9DKUcaAwhXnLZUXsnta3
NZaibk558yQQ8FqbeaJbQbO7m58j/BdTNy+O8Furyh4QHM4WcwuDPRTuIpGBQwj99mtfJTEO+jSv
gTebQd6DdKRe7p7BHA7kqRis3x7mw+jqzW4mlir7BllfwJpTULNH0K/Gc3O/L5Y22hixqmQdKXBX
bL8/SK5DVR9VxxSNT0VoSG77MJPDefZelp+kLWpmcqMhxlJYpKg0qLh2mvHKI1yq0ESu99+uGEJz
8yZi0p70t0ePbhPGlzDa0I/bkhGEuljbMgx6jRIl1Qi0PRuJqPwWJevLQlkXtKH2pv7NdaBJm1LR
Y+B3l0YyHqFPeqEZiZjW4YXk0tzf4fmH+FcoLCK2MYjKt3nVvbp6jOiOIn117fbo0CNO2WRzWQ1v
sCyKuYCXclCi1GnDHpw2fECOAy290vDv6XEPHCaxNy8vLcDcsd7sDcq7JxzckErVlsp3exddDLRU
fmSri+3954JU1dQmAeJVblK+DgJs9yUU1zqJ+IxvDwsYOBimoPIwDbQTH2DZFsvcdTk10ZjSzNtE
tbbb32MzBRXNSd4w+T5UsCZLoYi3gf7fvXuoXtFfEn5NkYfFKq+XhaPXF+8fWub6A5K3XuFVKcRL
nvxuN/PFU1IoZqU7tyHX9FzdiUao19D9Dzax2Klr/2n0ULlrYgtjAFnNXZulSSysG9MMEZBStihq
fpkYos5RuTLaZgHaLm3GlK1Tz1I5A4ECLoBQoPFGiQXytXdevWEf047n5vUv2dVKmTo2iMlgIvM9
b+efpwnAXmfvjrUkYEm65lbrjY+OhLFJczZqDmZciybXezOEWlIjLOm8SZqmM9HCSMgJI+xpfGsQ
+bkUMiun6EjBhVNzG6D3UAAWPRygvQtn19zx9PSsmMc6/+3531WLLIdJvXSeKaOIYLUw1DENtzQh
hGXHdA2fBh8NMhbjVB0I2+PmKhUhbIrw3HQoV5Q04kVSi25bUC+VmMmne+9apcamarrALJ74DbHt
u+W4pw7k2cHhNpanBVLRRp28dnH2oHd3kS0FDgdghRZgxn8WQBls3gwzMKsM1uBYZQiLGf7W5zLN
WEtU7CeESuGlunnwVHf2pYmPQtdWk3HPg0zJ/MiT43JVV+XzNm+JNsGvZVn7CXooJqGGqmvS1CKI
sEzAWfCTJjP+EFubdC4bM6GyU1iLDeRnLkExzP/t7CSXQPWmqVUhsOld4rmQApA/vCMa80VIsbNm
iKS9dLpf4dblA7qWHB6UHJ8oNNDsf0FgEhWaGjpWY0SLIh8K0gI2w+9EZls4LEoj4d0AFsoeWUA5
PPL7fLUA3I2wY4Xa2f8kTBTeHp/efk35fJnsURI0akwwEZ7PH5C7D2PzQPVP9kpVnOl0b4AasEnY
3oq0TFVZmYCO7A9VhJE38fmQr8oDgiLXkepal7BHB/pBGuql745/Uf0Ou4t+jZXS1yHefmqey6oo
LYKh8wWO0IU7Vr1/ijjQNFBWAG2QL0KjWJvNe71dcgy8Z3mP6IOo/zTgsiXrd/3+t806s/xfiJAO
/4dfT6/6bf5V9/LvS7esYRQJLs1VNr1rqadPEvFsTVUfpIjzpZT8lAVSil2XA1Mxs28dmSm8Xhfy
3WC5BsPsxK1XuRNB+JF5z5ap/BvPLT8i/xt1b/gcekwligl+Lyal/V1uyqsiBBWc5ypbseEmG5ur
Dl/izhys2FJHrRuv8PnK0PFlV0Jxbkv8JVgeTdEBS5f+HXXvBiJtwcEcBHQIVQucf8eWkNsiBLNG
xXUxpfjloiJGYqGzEuuJOVeJBkDdytA68ZxVK+39ZVOH9bQDeCLxthgujvSo44sPzH/3miE7mTNN
UAdRCfd462wZY4rZhRvEPXRyL7Kmx5MjKnXpKH6ge6h8pTZEIChe6yqClN7pBqyzFVM6QgVCMjFu
sseEtSTnmRicTIHmEIgU5+vILKIXKojIF+rl/R1o9dUCoheksx2s80uSikJSrsjIs9DJWsdcwttA
e6aBglmfXs8g19YuRlw+Uz42lRsFBKfI4uUpa+B+gA+y/99/RTV7JDirSLM1XFK0f2xSWEU0oM3z
PbUGyqhwRaMPuVhYrKrTSHnhUSQYPYhvj2SroI5DzCE3W2TcEpGTAWpjGRL5sxttZ5Oa7chwSKW3
5+yc3+Pn5mGPh0OswCN9SFQVH5lvhqO/N17fGeIbNMLrmxXptiLc9wcSRu/Ukxe44RoXtLx4zh2Z
iNq47r1gp8jBg0AgId9vEzgTLOMw8YNh4L8nGPSUH4i3DpbPlJpJDxJj8qCuw6tThrLX2IYFCTyS
BfxLsD+hEV1v3PCpodukShGa5ftD4hISZuDzaNpJtEBfEtyVL6pbUvNeS2Yq+H/Vbzv+m2Q2qQhs
H/5+6a3YvOl013Kx2razmVuCT8vR/Bpd9mNQD5/t5HFu+ppHJufHRkDnXy4mPE6juw0tHT+oJuw8
OGhkSBcYNy4YkJej/NUN5Is0HPq5BeV1/0OH0115v4tNo/4Np41RAxMB45kMN/2GEgi+W+bl32bJ
QYWWkdPPSw8TVPSYWoYqAYY5m7fQY5fIeQT2wPPvwmKFqLemhetqvP5JbLcsTND2uJGLkzncGZ1v
cmIO/k7Iqo3smcShKJb3WP0Vt9s/YsvOrm4gqnCVYhUbbookLGQJzu+LRbS/LAl4xxe6wqmY2gU0
Gv2C7sxT2SXFk0pchTXLI9EeVQGcLsLRWnsNqCMUpppQRsoDnrSVO6k4+DW+vbo6gD5f5gPcUhaD
C0p0rpoQjH45AHu0JzLScto2T5a6JuqwYg3RaeuR1xSZeFtp/t9wRSldKOM+ePPVl/CQMTWut+WH
RE/whfm9pZ1OE/KNZlvFtUfgUZG8/Hle7SQ5fLsYAkH8qHsUOPLeP2RtWruXxUGl0CHZDveXsxDi
JGyNHVMGHWhe6FVBEjiI9KegnIPcpXgIF5S2iKP1OuPt1u/FjF6hcntp5P9Ok/GX8R1uuQD9JOoY
OwMsqaI+kg5itPLdW8I1aimaRMgewxo6SpFHvcyqjbR5gEmJkRR3BlSpV3Z8+1Sz/j+T+AlwK4M5
BaX93IpQtuQ0z+8zJk1bCmO/eVwfzlxeCsANK3YjZXYAyBJOuau6BrwYTCXBL/EF7U4eCsiaet7f
HoAKGtMUpQJNTq+f1CPbRKWGanT2rieyLnqPhJiGTonWjUf7py5id72LvdG02Itplg1biikZu9QM
ZKJ5YWEdc/jMSX6rEklTfCBjeDXFaUb+1ic15NXB2TRia+vRl0i1s8B3Zpo6yU7IrfolOWXxiRGg
dz5oUE/Q95beSlQrzdsV4WOjAMSr6WX5vennxWttfqfZiG4/3jNFB11QO+Gb8PYua8jpI8Nk7jbh
uqNfCn2GWBpqxYGkXBA2mGF8MLRzRytxUUMp5uzGgKwHKRCNad8pXuOkVJCBP68hYS4L9uVMlaVK
aGieLACN5K4pSke/Jrhpxl6CgCY7eTmFSDpJIqJrC35FKgTegFJr43V3A3QxbktCM9sMoy15ievG
Y9N2R3mDkUjp7N/5C4PVqHkDmTyswaEAG9XarzAPa2P0sQ9uLkma5pC5QcHMLHLY3AbRVVAfM0Qc
KHNP4CHb3+hYVwfREw++1yRqwoGckiElfiJduwkkf+3wxXm+YSVLifZq8RVLf4DYywqE4idnVH/2
RsUOo+HBipJmJTSfiVTdGm8S1Wo95cRExLBxX28YHsOKeS7CHHsm12l3/D8eVcbLCH0Mpr8JUNMi
9l49oiwbsiHBN/kan8AGzH83ReDObNMKEfwIefWptAq+h4CLOXhxvjVGE6rIA67DbArTYJWFgzbW
+wPsn4+RB4hklEHdS1fuA64Li/xanj9WT/xR4P/I4wvrY5O2qFyVDoQep4B5Rd1YqNgwhfWYOxWk
OUfsQ+cyA2U4nY1KcUSMBZAcv8JlY+vXhVSHBAofSfLMJCia0rW0Ia0NX/VAkZeYPhR3RiglPcvI
RHZ8g8Uo7YA8o+GcJjNlaCUIv9IXhIq+z9JlNyk0YP+vW5IXwvSgr2+8W75IM/B+4kk4huolJId2
TEOYcLtzsOdhRDx2epnJfmLorFah1v2+DVMFeh+S0uUOkL81X0Jnu31uTBJC61h71s3ppXOTPemw
3JfyDit+U9HlwYyq8weHc8zHdB8Maj1u5SKD46qGsJ/eBXUSAwrC/wnark1fSpXKY0oCHxQxVKf6
RvdKpM6JyCD4RYl9ZXDL9DnXV8LT0rsrf6h3+zZEoDIiiykgwPofjTr0h2pY4UnqvgfUcpoGRQJ+
47wegEjMNXqeY57x/XtSmCuadva84kmsKSP7hhpO8ouw5QaPC24Ke5iv6kuwOnPz7s/4Inm0gJvo
7sB9QbTU/RsPKfudoTXu2Apu5VJCfa/RWhEy3QdLyT1TaJ3OTSK5FBm6MYc1Xpyz8RV9u1hDRFCF
WNjC6CADmMAZ8bMczbbUrdLZITcpzia6e0N7tzdZ5DidIbQDoia68WX+u+X1fzPEp/W2Uy3bNanr
rvJtnqmf8mEDSAk16wTol/4dhH/RYskdIQAGzMf7YZuDvx1URKCrbeZrp5A8SSrbkpmBBv1DhXMz
51LI+oYqHDtC/Pp7BK7lRx70wiDXFwH2ZPfiZrJ1PWOIVZue07w6zJx+04dqF8DH4ZQ5BLmOkbc3
Q6MV7lJy6nFEayo+kGgJ+wcI51kuf33WXflJofHN3gwMnaG1sCN62U4tHVbcF7ZZWhzCTMrQrnDz
gWAdzQ9vqi2YBya4vnEHXyVq5wG2nCHmwRTSps95qquSi1bnOwiOLv/P7fZF4gMAylh2kR10UaBR
aItHcVgmWD/Zp3jWKLUUnEHcRxfIUDydG8mSsV8eigJCaDk7YkIys1jjtdmjUgTOlZ+/ngJbhEyf
wxg0narnDezoPFWnhDuL3oxf4vYRzgeSaY0ibNLwLY1EObfAcafdivYzk2bfkZcB4Mh6hr/g6IC1
isJ6U0tiLhzjGIaUZydv11EP+Wi719So5MUvZX8MPyHLjvY1ssMz6LXNNPEUwXOlNs21otkZcQ9g
3I+Ysf5B9Q27bCy7dpDWAx2uE0uVQZW7mRK6A/lrJs5mg4M+m6xD1vocGfdTdxeo0SfLq8dKOsHA
scM6yaCUrm8cnqzi294xK6/H8mB4nSxIVFm+luVsSZlW34einSvtNEgPbJBb2MPC4iS/avCnlYAH
AKh5sIGH4rh76ln402zw/UK8/e/lTZbdVMC+I1Rpya9Vfs3ULvN8cf4YTeFjnn2MKFDXtQNFT+rN
3TvP5Zq8xFNVdbRTWRRVH1qFo6pQiFQYZr3Li0BQvXNAKRfNtVikzUKWC9ekRXWUEEL11DHifwvl
wnqSADKk40AhU/N4zcc2iVujzWYzCweuhuUMx8s5K2kdm+eyYmYv4eQH5SQLk51ZQ8fzUmpxqpG/
QTzxpXsU9yWs2jBk3czLKZsIsKxF+zqwu/Q0iaOJ0rPkk1MpGPwLxk1dcyiY8l1zu/fWNu0KMflt
xj0eHMQiPWzVr1BQm/BPo/a2IeTPkqkhBV9EcKrZfQ/efk05VvhWE0wNgu4Ts0Vo0oa2aGdUYr+3
9RDKERFvLj33HSETR7LmKCfg3mQPbSLXE+++3Om824APOrgZ2QhOeJzhh27y4Yn0Q/Dz6zGNZ3Ca
62bBATPKr4s3ZrLaVZBRoqmz1uNM/Zv0eg5zqn9WaF0lescHHMkAsAePHvZ0cBpleRCZR0Cj2BEG
7Sm7gDs82pjTnqcwFqqf+sFkakJL7A/5ko6E6UobVOMYNO9e1RWAgtS9eLncqrbYQamjRcDy3WOF
sPM5xscKanPJXUKOJg/+hnE87tsEo1B2f1M+Al/AI2jOcIT/4XUdn8NCQyBG/nCjw5J13wrhj3nf
I9GtQjfQQIFJnp/BibiYZmbpeJw2+nChd3FxUaCGsVrBJE3Fhk0lxCNkg6ujPmQ9RV2CwUcWU0LQ
hIH0x8iHGFAaFRniF8jbbVaMbtd943wJZcVJE4li+fjlGcaDqwDCIfKRxsYjqM1+AFev2gteLx5b
ZU/fTCZl61Oe8FB+M37Mvilp7LQy9Pngpc+14BZCDf24H68jHqp1YHLKShugnX1CiGilkB5FzE8C
pGcyANR5fSmUjf+NmtVO1XIW/O5u6iM6aiYivL/pPRCBxX2AbuERZSS3KCtoPHIghhdqLcZCY+bm
x/vMgL9a5pcd//v6j/fEJ7ZkwoBaOKjeciA3my57n3tQgZ7GmC2mjQXM31V82pwSQmJdPRO5cwTf
8+NQItJBE0JlXGtq3Oyy2wiOqfZY/PE4qf1HoM53cDGpQ39kAZdEQB0IknMBBT7xhM8qLpsypLRo
RlGj39bEuCmwcGmq4CVT7MPIXsS6fHvWud61+3sJiNdun38xV5iFvKpHG1Ugxea2wlfNaRRYG7A3
NkJmNX5nIp3X5/uxs7CC05P04Y+V+w68Xc8Vrqc7GdLxEaGsBWn7vo43Tb7wKyQx46oVUCyNEjlb
FSHYy7Zr6XRYWXfeY7dd9AtyiuP5/wTshR3N9/jCPDTLB04i9N3e+ipFxbuHgOBhZLh1gcFOKbYM
clld3szDnJe35S6iV/ZoZE69i8sW2/mEudPC8Eme/9+Dv/93COc3+MhmzVLqTrxcNzDRYCqCyesp
nFgdRdMRRIr7LQtwROrcqhbI5uXaHet4JEKep9vMykUxGWI21Gch4IraOgh5Ek/3eNIEMIX+uZVL
dBx0gCq45m2Si1CVX5d6H/TDnikO+oKRvJPwsHd2LeVIwqXKKliAvn8nIy1NugbZeZyd18cFJbKW
1kJDagqjl9czYyIRes4C5ZNq/cbcGnxTv2tAe8SEoblmyUdV4oleeAoQkOqwr6UsKrUL0Gj4pSMn
lvouWia8wW/FwKZLoobKuYvepGBK4Iv5IaGnMGVkDV8Hsw/yocp4MO1F8QOJy1urZoSF+4MSEfJc
x+QRTD8dSmwlEc8Fh7pWRUPhQ/sF+5VvSMiot0VRGzLwCoJejnxIV2NWVgIwoaNKONClz3rTn40V
0bXLT+hiXyGKQDKpBNYz1CWzXf0Xy6OiQaj4buAzntUdbs2Y/SIXFHuxJZuOEcX2+35YKHZqkR/s
VqNKVhl8deyy5Ee7WhGkNcB2wnZMqTlX9bKy1QyQXOEhxCHXbad3ZDfufILR2FDTY8OY/uFcjy6r
el9AgqiPvQEbsKQEwY9i3zebpuT/deTYYYzdcfIIIMcGaq/iImEJHPWfZ9Yij+nmrIdmv7LWdidG
oBFq0pUYt8ILw9tsKUpQyrEmpzqbYVkOGSZHS6dV1+kgxdR2IodVs9h3tBIBDnXCSFIccC+MOtDd
P7zGCETii2nQZpYWYia9BkZ0xDWUhbg/Gkh5D8MlKE+tS+5M//asWcAtFhdmCmxLA414jjpPWMF+
Qz48xS0Fd407DrRdzpV3cRm4jEJCdvTPFdFUAzISU4mEjK14VYa+YZW80AaQrM57AItT+piNbsdq
rVWwyiGh8oPqY0eVP+YgzYpAXDbo1cNIBC7fJNHaxPjC0XKjRhFzTWbpb4E2txBl7zwQK0CTV3Av
t1adNCyAPqGY1JDKbcq1nFXfdG/Bylw20+G4jMfNQD8gRlwB63aK9Ku+dnVElV04cI9tcXhaxq/Q
llHdKgsf9W0RnzR9v1hZYdLnUiQE4Ru/4ajMYq7F9WtVOeJc8TV3rzB/DhKOOypOO4i+3bthKrIg
TmpP+Yid/YAGMmpc+T1EHUd3MMx93fkn2/tIY75SNzWmLCiG0U8pW4fA8d8/bNfjID2Rfl4b74WK
lYfSFcbU1Y+kuPVlAAKq7wt7SzTzqc6AbddCSOhonOkz1cXLrQGNwD4Xw/TprvCVO/cJ/NcVdBcQ
enzr/+tAaaRrr7MDqkbO10I627SliRtTTElbosgbgKKFTSH2cgzezWOnTMER9w2IzC90MLUiSuZd
6W54w7s9eN+uKIqMkJKZijtXDYPPO1qswfoI6cpsJy4eN2niFp+z/2hOWjnwOKrGJigUL9NRd+YW
GCiA9t6PY+d6bNxXjWjEzTwQ84/eaiKUH4BERx5RZTt0xKQIa1GWePeuB62sv9lrnfGNjGgDfKTf
ksZcqurj88mGXnCif9WbLdSRdNWxGneaTdcu2hLYjZpHEh/Ftg+owlrBe0tdO2+MG0pj5wM82GFA
APVvff+qKIsVJgMfONxE5Q0uozCUxj5aqz0LKpx4wsdH8ks87K07gnExm6AD84pRKbt4cLX56OmA
E6pgKBhYdk6ehlXBccXI/LnyUdiWUIPqzmrSl66CCMCn8jPWhxL85xsRcXRLiuKddw+wvEyTGWJX
ML75dC4Ih3emaC5Q2/JsacF/DCLTLKOHh6saD7KOuJBWAC4YrcHV/EmEYhhv4wMMVqtO8FdBD+EZ
dOLVuuSLbquA2VyoDJeJquoD5EHCSVFVnvS4VqW0ldnlsyGOXB+XCsfVbATfwlH8YfjCoIx5o+FC
BW0GVj4Z89cErK1UcSlBrhgvYIZuO8U+U7kFvLQ84K9CxtHhKfBhimcuKzCzcSLibj5sz3/b+9Qt
Z9sF7GpjgR0akpJF6wuSiWnPngcjNFqCV6Lb9aorVUse125yN8K7eZOnMT+9OTPZTnd6Ch4CW1Ll
qkbsCaMiTZrF0d/w/xacUt3cusyE0nJrrApW7ySADeL1GJ/xAoW506ePql6HV9xikH6bJqoOzgLh
A5p2ZwqmmslxrD16wVHfA8os46E2kFBEs1nix4vwKHa+RcES4sIpDSlwKIH8uIw57U1ifOpuBCX6
0EkiaGCMaN2tciOpemkD+36MHulRRvzsJ1griOIr2LeOBePdsiIbxqLHODb3/+/8GEydRErbfS2I
PW56AHiu69MhQ7Bz+SyqyOHeKm2jcwZuBXd4YUFyfVx1dIhvR/MtYa0hCE4spy3dFmQSbpJEgGUe
mfN0YP2UuFI/lppB6SG0EHf9ns7MHLeQ24JsjEu3lvvlYjY0MggphClU4MbHVdMHzwyM8P3Mm+39
TyzoUJ26u5GNoQSQ7OC2QpUJ0egAWh6fnGWFauqg7kyOP+p91zp7uj5cUlwJPzzvdP18eCQ5H5kg
yVePpOBW3h/bAtQzjxRh43xhvDGUZtSQjpDuHCVnfTS3nZEYK213M4xfO69lSJQ0US15xSysKXzx
j5r5cSs0wdd+Hfm4G9JxRzbM9kC0Rc0P5XdZ5XPONda2BREXufGxjnujPBCy3ZRYOPoB7SlA03F2
ZO0RDQuawb2EYqs1UGsjPpBsVzYGHAld3R2PKkT9L1yM91ssIz0uCRmnY2/Qm/aQnr7bz9qdaPwj
5Ueunqm+FpFwZyHru7SacMEY7kRQ4Ts1oquY+M97qIdB4BtDES0HG0yERqt/pTlrMBpoQFyXNhE7
EBhaI9P+vxl8IK2zlqSWu3GJaVbdpLx9vg6rWgAEsy+agZLEyc/pKpbSrmhiP1iUHrRfk6JsBYk5
JJKyTHKVj+UW2wssj0uppgI6dHMiM6LtMdoIMJY2zp++4YZhCQp+dRCKQrhex8VObKwprVc/HdfP
WKcYTCVxjWK6OrlGNC53FqKQNVqtgvK8/oMD8G2p3oMs+ed8LVaePcbtvlWlTP+UrWwgkskEm4x7
4Y6TlmQRP/zKDJCV71QLq52mUnfE11ePH9IyxDj9dXDfBCFLJX9DKbBueGiiVsLKEb53DDL76xZ3
dDfev5bh6h7Jpq3LfqrBPkrO5hXkDTG1l59CRwJ6iIHYi5eJeloGo8lREoPcnNEhPc4j6zTokaGz
3S3aW2qM3qgdQAdk58k+XyMuJFS43pqKrDo5vMmPH+pjUwT3RalDkKVrtueT3gLvnHkeVmFOyehh
gsRcgBNSNp21eQP2/QC5hLb7cYtpDeiCcYr3DsFWi25PkpI0Meapzy9N3/Qh9CTAWwiZalrxFnY7
JryEPQVndgYKPqAo50riaV7j/RZinEt9jiuj7TL2ofifbmL3Gtm2MuFgJSxqtZYsYnGNS8hwPepv
1kF183EE3rQjxZeO0zJluIkpBI6Aq5YjuAoUo3DgdBEn2Wa1Q/rlmDNPjuYAF8D9yOrny2SwXHLa
5e15V3RMoQKr1ZX6J6byIH8njlm8yFJ1ZTuXmVKmLhmWbRi4rB/cwxR3aEema+TKVZ7Uup2OeURH
zr2raeyX5F2xp0RxQj2uzlYUmE0CZhPrLj+kEGYWvp3IwHiQ3dHS3PwSAkHZMBwQ7sHALCxMy7io
hopFWV+S+7MV+hj/g2d4IAqJwROtZWW3eZeqOorIBz9LNUEBcj294JW0P4WSa6HjAgUKBZkoqJHf
BpdHsXG4YCXPDVo53oSUqaP7ixPmRZKnr5wF5rVpdpLneREMfKURG3/bp+MUDVkLpz75ylmS/NAz
UWgQ3dO85l1eVDsAO/aXymRdohm2BBsSHKmlguhVtIkvE0mMsTYWQ5F+a3f6OUIb8AA0ro1t9KDq
4XZh6Sclo87QkbUV9xy4QViKdk0xkWEt7SN81luconipr4SRcahXFDqoxGuAxB5DqQaUBn6a10hZ
N+/mJJzs7R1rGuNlS2MkkHM0BIzO4Ha2XrjO/o2hI1JAyz6Bt8gXUfXwSpr2Qy4RdFwckhqgAGg4
fhiro2hjmWNvBt8Vk8aZsUW36BpUxgeEu1DSC7mxUvVVqVQ0P6IhC7oOBc5BEGZ/dIW9242sKz5P
+2cUFV5HEXgDqLYZZFbHx5dXkX5clJMBSowA/oRZ4mJ+IWNRGwXnmFFkQHKx0VbzCION5VcvfuM/
+AB9s4kvYG6Cbep9v8sCWsYUKW7QMvJwTMeBiy0yh9eIx06qs6ghlKcYGvh+mgs6o/hQ7aUY/JEx
C12yd746ktO+HqobBkmb3XCIPRIMeFXPpW3QaIN8FUvLlRu3Y+Gz+19iV+BK0ZJdhiYshce+gOSP
+c5ap54rDkcRRztmLQDwzVzRi3/kJZVHIbhfIdxpzz5jCAjlZeD50CkDbvlFP5fjsA1Af9VKWfT3
OHkD6yypVMVtg1aVwZtjek+qDRM3igrLo8sCR57Zp5NXaKQFdh16ZNtpoYdHmFxTf3iukjFCoTSN
FdEJAdD2eHsBMSa8NLf8KQcvDZ7LFXxCViBdmZ5IPL+8ffVR4tbcU0PrTgRvy9Fn7Mk9jmOF7BHO
uthHXElCvCJo0R9brF3Ety7WzIjHKM89rtw09NUj8T9G9vPLo8zPbostutKqHbx9x8D1H/LHj5tA
h3MTtWY4YajHC6ZWoz2f6+1zp6YoTU/m1895NJZTIp5Tk2bNiPkYo3wnvxDBz+kFZLT9QHtURYmC
bWn2qfr0IglbthP3CNEzd5k02r2d2e0P8dbUlaAMqdz71tUaeob+zmrxicTfvzt2291MqSIomtpi
/gaqm/pB6Tl7p7swJ14diAMXK6FUOd8Ik9eG9f62FNqnCwDkXo+nggQEDF2EZJb3kysXIIurN2wP
6tpuHBI8q4+yhQ+2WI9eSkWt3LW3XtlZ2Ip4O1TC/jarHHkabCGUIu0lnVAd8Vof+g5+xWshEojW
zkXW18Kzcjd6L68jYQCuITk/j2paMf2T9Z6r+GeeqNYmbjIqybvBTVaziR6czoAkGBTibw/IAlES
SbT+g+0v0oLbKXSmtZrxmE8X2hBMeJSbGzpIYmSTXOSqTJimo654MQZuHqrjzAKcGfKhnz1Glgyu
jRj4AjTCVrj7OwL4rWdX9cSgG/P7mIUJwQN7ihX+TzlA+Jkps4OaDKI0epmQspPUsy39OGFF9XOa
AV2zigPzGCvsOZ53nnnsfEMNV48mBSmwi5VFppTAizUuk8VXDmZMS66SiWXyBx0fI1ITHOyvB6Jq
qPOiToePrw/rLK8wecQNZ8S9Eh8lnr9KHjzCZ3YtRgZxye+fplUrCPIB5lysZT7XpYLfxeiN0+vv
iZXLa4DdCmbamcU+HbudbWlOoxcGSEqSWRyFz0Yj0u48xe7LcKOXtT38lmO7CBxYwRN7M08eFu+d
l8Iw2/ve2rdeY0BYdV4HBQJsAD3NbtF2LPrfER3HpZCZV+mFDcmSYavzQ3ZdH5iPsrGL310xthBE
PRZU0USO+UmENmCgnG8Jg3QsMDczlKBEPmg2I18vb3pd0pipRooU4wRgsvM79YtZqWC6dsw5jCIk
nvFJFNl1ZzYVYAbs/A6pUL5KgoN3wmcf443rzozuaF+rnYMtuZ588A/KwSjOjpEQXrpjoOUQ45nx
ODAdirFjsd/3g3Qa4Ln4obAexsB4pKrQOwTZ4inHfFnTVs026ltRdntT7HAJXTY0tK3wTU+Xlc80
+b1Sa8SUElP+LR2RnNilymDspOO1vGa5NKjUrMclgBCQGha8qp/N6IDxhxEbu7mcfbcI43ILX5U1
2ceqjmdWwgM2VqPivw510TO7RRBMlyK1B39bPrjLjoRtYBsUhkFeVmITFxTnQ9ueIQ1Ci3R5Uz8n
aCPCeCITeax8xe7DwSO7KpbqbJ6brSQpyGIN0FIEfPz02ZUFNHQ1irDQlr2TC3kR153afKtJKPWH
sXm/it4fkEa9tzbCK20KP7Iuel3EpMbq5d5pLQaZ70DcntQEWis5btyI/w4yXyYo3dEFpgMvALlP
7kCyukQq7Msu11MoSo+5LSxYFUKdJzAW9x4iPIxXHqMaHmY7aTDff7TdorOXp8G6mkVhuY7dwh/A
Fk1B+JdA9GYQXZ/QS3bou6At4CBbuoPVon48v2tiM1dq0Ier4cjkR6Hzk3T5uNj4PKNNIvsYW6Bb
p//DoGy+7JLnb5Vn7ui0kAZFfgElvGGqNu6aa0jHeQ+RCjw2vp6ioMSDUgb6Fcyz3WIsBtZ9aLqc
LsXVIKNbH9punJoAvXOM1mi9gjW6Gk9D3PQeyIrLd/1Mk+icRNcUfpGXwIbswphpLgehe8u0Awtt
42KldQcfMNKpaJNZn12t78VoSJJvROtbCehgA5J3nL6D+ylJ1eQtYKeb/TN3LVuujGe5Y/rew00G
DuvyXg96Lfy14H09uWyV5RujKZY/cB9ofrxhrvpclMO6uf6Y9nVlXNa1Zqpa61oigdSbLqlmkdKt
Z7yyBbO+4KPTtraVEe/VHHBDvNt3nI/uyf9EL0/qXQQ9i7BCoRv6Q0NKhTwJOeMq+SZPW+tbfrpi
twqGXJfOJCuHS0fIRaqI4xwPz/mQ9gkRbOACHTpK4cocQflZtD/9QIa19hmxW4Xyt6LlkRUB3OQ5
glDpFDwVyXg8FSDUgRNnoqUgUpVABGmTzUoamtM0P1aGnUrMr8iArjC0rHou3rzYmrpusoYxHKMa
HGZVTJNV4lwnmrWlAH+7llLXygNcBPu5sikn3JW8IrgEUX2yQwQpIcqXH5IHIff/RlKmTD5v+9az
gguKqDnQnYwboqujde+VYLfSddn6QmSemvrViNXRiaE8txOQW1UFNKW+KEBqU1D5e7ScQWZQyoiY
fU4cVHpBA1cCB/Q0fW6Tj6BBGQPAy8b+YsN+LLhE+WDmaTphpQpOinOEbB0DOzdGN9wRQTDBZBWs
yB898p9BRw8nwpWGOLoNmN1fcdiov6BBz7NNYZ4Fus1m7Qx+RFdvRsNDVSyorK4f2+zyFA55kssm
mDOFKSYKveSAzoPzJgGmoyqKlSclUsXC8YeejYriYS8eH0NFBTa0Vt6Lqs7jqiBXb2JLoVF0Cl0o
qc/T4HFjTx0QFUe6Bob5ZVV108Oj2Z3w78D7+LZ6PFHF5k+Ffs8m0fpixEudmALVffHJguOW3cKd
uyEZqTgLqdfG+fb1+GC/VYG16Vm1dU+fuR0ck7UB8MFskO4sPVLpOj0iIG7rcRFREgDURbeb/S7t
PYHs66SNhaPfnjGVpvpkSV+kAPH0Coja+LKoSGEcY0BfeXGj2vtqbkLjIemMI6mExlStUjaAsMpv
jWFSS+KLVbhMGIo5QGZegucYd77/+s8YDwf+NB1XNXw4eR0zOKi6TTwrqsDU3Qx87LptXQj12GdE
bHK26u0mzyITNraxF/NxmSupW5zNirVk/8/EPCbJrBswQiKyU37HAWteOHi4BMYuFvS2c9czl94Y
mEK0RBwNjv4wBwFNCtoyH4HDHMRFdIqcSOU8ym1xqXyb6a+2/8Uho//NW8qobgInZizTN4exdqvf
i4h133PVD0OZ0g7wX9CO8Y+9hsxrQ+ySQkWQJGlvcn9OPWty/E2C0jeJesh7FrhLQ86gDJwdx6Yu
Pfz5Lt6APJiUadbKrYVH+OqRqD2kfO52FbUDxbjxkwYB3J5QlCdtYKI1KfTrqCfB3nbnZfHABw+R
Sehw93cJxazY8+Vi2eArvrfh2uUIkRohrzhjMYalEW7OGnYa4LUcZwYNeLgIi9ZfYR3q0+MmDCTQ
N9YP6i6nNpVTR+14ZgVw1dAMODQJ8pP//dLj+mwSFvgYUJh+c/B89nN9eaX8UB6ZvYT4g8iSqqQz
tkFeRCEOVQ0HoGiJmk2agc2MqtO688LjPSg4NHuF68sh6EwIrInUfc+OY64ZU3ZF0n5lJYA3G9dd
MRW2qyBqPzwqIxAXsdHuqBOhWq4oLW/qmmSaNpMscz+vzlI7Ingw7BOgFvJZwtiS1UUfmYbFY1ww
5LZ3R05DGPRpiSVe3ZvFxNZ1PiF9uNOOARhlE5OmjX1wFYGsJolbeg1uedvW5EVM7qYDbhLkwdi5
eE0Ijua67FIR3tEdmK7bFBMCRY+OkUTUi8nhOHEEPQbgJjljKESZP7/HX9ak0seQHPAqXoOJEYaj
AbE6pmqY9AisFmuNsVh1iFSYYQx7dkbNdOy8c5pQmX5CuvXA6AFXRFqMupxD9eROx4Nbj6pUxZ9G
spBdbQZFtprnEh4LKOMSVnWP6QNvbGZga6WMPElZzFhTTc58uJ7C21Iwo75uk7zm0hTfxegvyFXq
bKXehlhl3eZzACffynnS5VZ0SjrVNa0IsR2tvPHS4WUdkBXbJsj6YxA/Pw45Bju71r5QET6RpWsW
z+p8f8B3+9DWAmI8Yy0WUskRiLQh0+ew3l+yzQ9YpJhDZ3eOAiI/deLpH9hO2ymih0HbMAE+E3VG
lIjdvcABuqxLmvvj7Wm6PIhjSBhWRM3q1WtXvJiRUXG68UbtddAOw5z98klUZaCvSR+dT9P3vFJj
3gBiSSvg3CP8ugbDzFF6EelOUKTRL2941XgCjy3LnW5Ybp1ZCWpY5E5NXTZrT1skk600eAGfNu0A
WnJvzVn3hiqwfYouHcQX8s7KpnZiUR3iBjEmpE9pM1eJ9VxoseLa+NAzawhPAUBzAaTiit9AxX1J
cfAowqNI2sDtuixSddf1AvTFbzB6wmOZP5cw8nRKZ/rxlGUkOLwBCtR63eLVm8IQIvaX6hjt7jMF
BPaHVatcWrO8KPZhoVtSQWeMqxUQN8kiOw/cI1El1TW8khV58gImASnM2JhHzWjiB6cJUkBG0CWo
Y9NM8DQb9zHkO83S/16jGDydi2FmMjusksdVn92Sr53mFno0ca9CFNVEP8UJecWjDosMgpihjaob
s0IqbmM71Y+n7qOl5uMRQ99b2bzdB3cadzhYXwFZCx1pGtF9wliZJr82qL0rWC3giYrLpbZkizOm
lxuyBBRTMZjYIR7R5sDMphpS4xuKWGmgyww14uWtONFDmfPX8R7CojG0EPHR8c66adrI5ZX3hBnC
I5MF7Q1Oq7NIA/hL5qZp2nbsUUxWyszyZbmF8ZXBDVjQ1Whm4SYWMKHS4P9k8rRSvE1ajaKpqjsP
zORpEhcHk2RrjwtNiOZbUPk3Akxo7IAa/Widmg9ZsiumBfWjQINIYOQBB72lqtLqcOMP/EOlWPJ7
ML5FWCjQbEF6jXZgvzctk52N7zipH+956f3gPmq9Kd+BLBKvllqNTNFV2f/WFN0P2HX/cU1+n2tG
gOq2OvD6CtaHcGLY+bgBK9FPRitB0HdZkZ3XG6VEAH4VNul6yUCKjLns2TuJhbfn3O7z6o4ZAw6v
hSKncGlUO3PvRSfb7Up/O9HmOkCevo0yzwA2wXjlTRaTePkbHYWRZVcNQgvhK4U5/2qao6xZFOxk
UGTRnp48wCMuiVAlvwOnS+NNQBX3J8hZSzoIASOvzt3OLIKhGByB2TB6ekyp5A6zp6ixxS5mMx4O
IIMnLlQHdErNN3v+V/Le+I625FSP3BRdBiIv2gWW+oGfG05TgHYq+TNGvX+8oydlvg6iID9TjkdL
FvuHp86r9OgYIl+lxBzHfmEXYu1+aDg4mYccTvQqHoWBNUd84EAzXtHxRY9zUPzkrBNEms82J8G8
/XfWmByGFuXH8uRKz0tvUnn6BA4ix+J2lrlsj6Fn32J1Quo+wruTdMui8+y3sagEGRcigdgGMo+8
mEFfJEMjQ3ssz+sAXA/7U80QNsfJ9kNKKX/NqrwNixFGJKK3Nc2R18HnsIUE5yll3mvkG9PBLyL4
XRlFF7xPK3YJvyYT1mFUWhfVrbpsA5aPqEctFz1jkaDUlX1WItMNt3nb8TLRsKQ99EANXX6PzYMH
m/MSRkFaY/cacEslzADT9q2iZGT2KCrNyEsanAoeV6mHbEmnNZSjXcfcv4PvD4YcUjBte5XrBSAh
TnEVlxJ647hA996nGmqpHz7YQRCziOO3RKRtgYbGXIN/9gAA/Qr3XUKfvJBgpXj83pZ0N20sL3Vg
jzWWcQH/XeEBemumuFBg9wW4i572ylRJNMYwVnGX3J3wCiL8S1Y3DWLZZjzRrqS9Ei4mILB4traj
jDvWEGcTPUAUB5MrfC725P2QdmtbZFRBnayt+3kaLuw3ZwajenM5YZVQ1nofELfC8AJOnea+Nvc8
uP+oZ62IJIKp6OoqPbokUTEtlzErLoaM1oWtlbLy4z4sYgGPDXYIhka1m4afdGFgsIZ5bHtbaUUN
5b5SgzA176TFE42G/40MXsQEqVQFIJFaHtvaO9TSbzQlDKSb9k+jQ0x7KMfm1P7wAnnzrRYkaUxr
UOx5pPqGK42fBQVdbZJEkUnZAshJOv6ELGovSkcE2vDcgXJ3FtruJ91vQ+rs7arrjEqocKi6az73
MTswerCCYP+qdXs3pP5pUFTxoH3WrUwGJpxi75rET6O29ZO/3Y1gnTYKryV2ewNLGMuBCMEfhxs7
wmdLfBjkWVDOwP6ZNv1cr9FPaVfHbwKx7ZRhqSCIEJofn/4ej/OO4pzQXmQ3NaIbxvBkh0Bntyy5
d00uwd6rfDEPn2IHSLfG9NyVT9Fqb8a0eWsUQCz3C9BusBBchx8cLdnT9JXlRWe6IPhlhREC6zmN
0xPtdjwbmz77QkZnBr0yyfaKuvQHLExSHZruSbjnocYN9yZopguVSJ5sc1QD4EdWEWv6UyfAGsrT
8eHVBHO/xusjcjJXV5W797sujJmq06OpTQ9MkvgElCm6pmI3UstVLNfiUu3cpAJojs6dJwDAJ3jB
8IzeGd+9GAO9Rgot76dnbsN2dVhILtkufFA0jCYNcpJ6CMgLcfO0hWtaWoGUMrsClk4vz8sntC+y
y7h5d3UzxD8jTAGBoFrCH8dgGuNc2ry/7p8748plOWm5tG0Tjp6QC1qeEJhbWKxUmCDjLWAS3x0K
vHCESr8wUAQUmiuIFlIsFzVKQWHb4mSSux5U1zJz4TxaKfy63FAAO7fI8hr9ZBWjaPAG/lJDivkp
bjglpeCLfK/91JWhluHF9DIwmXZFSqBfT+gJ4prq/hrtOOK67dwY0ZJbD7m2f0K6ktsN96LChW6N
h70dRlfbrELXCbDi4H5S8VQ89kOGTNXfZ9qx8tu1MbDlxAuPOqYHXhzX9BP4mffsh7E3LkmW9cE/
YwoLZfQpMRxajw0H3UBeNgCott1T5t2jyUQ9NQIemEpjJrvqcxQcQ3p13fI7Mbab742ND7dku2gc
igwymmHdbz4Pe+8DF2rIQshkgFTS5S+CJUwzKFEhEjvpXTSX6f70/lmm8PtLC2Ahk9sDvlVmE/8U
Cb3O+ehuG4Iks8oaMACdMO6Je+fT5b1q1TGMVhB7BZkwRwnzY527JVG1Gge6Qv9sxbzp4BD7Ce3k
nobukRkRIYdD3QYPrjEvMcqoCHzK/eKfgLHsdS5bn3uFoAyyOd04S3sjWQyLFEMXN8/asUciJLEE
hLjy8kChEXUqf+2NMD+M4TlZVCbnuA3RqcZPZ4mUkKcGaY9oJSn9ftR75Ztpt5bAxdOY7Jcnm6zz
DwcARVUPvv7cBr+FFagyx8BZ65RSKbt2SiVsVRvoY/4zukxE5PKjgWjC5S58kSJ3sf+4g+QUO772
zrZGG7W9g9eSBpKBLWpVSyc0qa9DbzfZ7nW2TNQ+0MhiKOfQvYAUZkYqSZNUVm/IXsf4RdeK05yc
VtojU7pHG+y7GBh7YOVZTxZDWVJrJuQ8G7x8XlVujEUuW8gFEQjXgbtw9eMppDthFqyScRi4wViZ
SOYLK1GU1ZX6WypI0/UJZHmKB9ezPybDg6Jl+YkhjXZS75bTU9mjePRgS7yNkf8EkWNuS8gKo2zx
5iLKbBCUQiILxTh1LOy3uDxAWZxp9yjDTrD1gK9WaHqTNcc2eHrYiBzD0ovb/4hPWKDLapwOquov
GAQ0anYsJcaV7v6ELe3LyVuG0i9Qh12uvlnBhpZSV7LqQIk3pqdyWCzAEP8NLKr6gpaeFk2cvlpv
TSbCDk1eOYt0b2QjRIgcrgc3NcYmEzvLxwLLgV5DliOtN2vD+Q62BK+Fb5tSbw0KlArwbaXn+bL/
xnGOiRwQWX2WwG02f6nHYjZkmokRxv74v10cC/R5mblwdWTThsI64c6D2gIKjEpp3Ta8BTqH1HBm
VAo70W+zu1f/UOrR56YVEr5CsOPGyYfndK7Qgl9bZm88Pf2ykyMJWbHaay7zqFh3qBSkrD8qI+g0
ykRh1NPmqcvPe7SodEilW6fd5wCeVFCn+ZYsYqP9rAFKec3AWOElShDiFcxq94yxnhfnaZVqb+YL
rxIFXXHo20x8ImBxZJ/2jD6/4SJ8nk9a56L0Ec4olTM64rHUkD4uqBwUdbHzrci693Q8oFesNGEB
LoyNKEc+S7Ua9Pq9cf928W7UkbOKWwS2cp0cKZX3LPIuBmtOjUgy2NGBeruZyLesGJHDzR/DSGyu
CRbTK+Ll++B2MO3gKbJ6Z2Dyspov0f9fGqdYkPQUCu1pxzS0bkEWXINFofpbi+a/HCUQjHGTcXaI
6BC74ZXullFlokmSAjYRFLixIVFwyE21G1qyL4k2AXBzAgJNLTtE+sJMO1CIHwQWlLD2z6k67v/o
YAlaIP0mv3XH+kGduT5HHjJomHTPt6qyc7tUQJueWeyVCuHoHH+9suYk1WVBgVKepqfehzSHCc4D
dv3rtrrzfBy+AvkpiaudT/wI+hRx7SkgdwO8n0CfTpVTUcwQ3ezxC+NDWfnuADpmJeuXWC+tsN/W
xMPKxl4a5uXqj7PpPZEgvuyR6JsJirfkxAaoislwdoytwU/8l8rdFBQkkcp2KaeK1BPTd5SQPG5e
KR28irYSIjEtiBdZi8MZucdRxFJEgBIzOH3VzEpBohKUALst0MuBcdP6kCIKZVBM8pLi2OdEdwCa
nuqJ3MWIlq2uxbkKDcGD/2oAF+XJRzX6bXQn/2bk9vOKy1/f4dQ2PFUrYnL/vFzZpZO2T9YA+OY2
Ls8u4EShAXaKttnDgV4V+Kc5wy4mqdooOd8BNxnshvfeEEoQllwC9kEzqxGrTK++95xsXUdKySXc
vRqyUYYz4MNCkbYnYcHOTGA6uvnChoDpmtFAyLK+ylkDpotFOu2USTJgrTdk3mFnQsWXMrVBVUGQ
gq3A9ElrbVjlyOKTrsZNcy/jcvB2UAsMUTaJxyg+M971DIDpvmuDmIxHASV1P743D1TKxYSkypSj
aCebQI3QyZjxXiIkzjGad5gD0oj59a1cOfiiW410Id1UYCjX8fEq3cEzN6IhDNM+WuC6HekcPM9T
X7N/HWZYn2Er/o7e5s7VmX7IKnOiwFgQWzO5bPtyT/Skcj+Li6LK07nQ+eaG5UKMDA8zz2IAOZXe
k7Ouf1KqkRVxUWCzZ7hCPs8fWmH+VZtLQGbB09DQAH2TgrrdqkUaDJUCZ/bVqrgzlmltCKvRx+8A
b6MzVzpGONmEKW2QJQUpsxOsRZFEjgRPl2ChTcoKrSUOzDPrZojeBVsWl6Z4vPiO8/qVNrIjnm7O
XAnJsYEEGZ/Axvllt7jV6aMkVL9KXTUdA0nuzC1QLzHocm+Jcyd68Y+ZugJwdLVnoCK96Gn8MjNi
v5itOnQyGdonDkRQnKVVu7e+t1QPuKO8ykv9XjUZJu8FltirmoA6lWPxBNAZwV4WS3BAFu/Cxcxq
OENZ2rU7za99/siv96dCVaIcxiQkCIb5s1AsOnOv4uYaqwyoUQDjBUp7ER6WPfXWGIxaGxVok/Wm
2uv8Nfw/QN5EGubO43OvTlrgZJ97EsPndeJjrJsXpNhg0MwJjm2uaj9G6aXTC/5cXaGknzAbVYZY
k9bZ96rYQp2f4jXTzwxaDozW2HkPz3OTqy8yOc5BHsTAs4LokjAg3cROIVUEqwX9XfmcEb69Uiec
HMRQrnodcLqXbVDZ3vRSLMQQXzT8T1mKOqpQ7lXYK6G761Rp5oymH4G34k2csE5g3PoCWs5Zey02
qstkpiZRwJJKLPuB1gd8xlpTZ8kUGV51fLCuBgXPMRsyyexQXSSif+rGEqJtBZEK/okYrry/whkY
oVx7HXOE10zZgZVfGeDi7hHnEmSshYCGbMVtL0Zn0RSMbB1rBbF7j1UjGFP86i21e/Z2qY6hI6MC
6LzlJnZwZU894Is9E5I5v++fGHlBM8SFjh5D/SP+Wu97JPgxEdJIGQOunpFsZY/pFRiLN4etswM0
FKmt/qQAZjtHQE3Zb4hAuKx7PNQB/6nZGOwXHF4Dl2No6SL80vx6Q7Azy8qj9xxHXQcavARkFdHm
S1SzB9M16OK9u+aQXjmElC1Ehr5IEGtJhJsJXYgO9wj+eHl/1bYKg67wG0j9qKgtE3rpq+VWQ8/Q
DfyrUj58Az8b8XODDN427u+JCV5V+giUTTN8T1mvCowI6TU9Zyjd0GMTRq80aWyA4JRJ3w0K1qyh
sIf8ChulyKtfpM4qh7x1MPM7UhR4TN4iTPsl7iwaNh6TiohAd0StWj6eJPNv45TL54PLbktbV+Hx
kRwk972qEb2ng6VK6IGRHTHr87iFpdWTVYqhMMyp8RFcfifvGxNG3Mw/Sz97IoBLQfhLUwJl8+PW
To39DHPOXuXpsq87w7gLEmH/N9MvDjXM0aEpwSuOdypu7/x37gZFsxvrQJgMJk9LH/XcSLqrL1Vs
p6aRDPgBnyc2uBebkobUcA2p/kHtHtGugrALbMWNZ7cF1tSSuc9i6cUgGY5/HW8rOwS/czv9sHcR
LtAYL0Vqz2GqP9Tdefbc9J2J1yFMbP24//sQv9wDAO0iyhIPVHy9ZkV+NSD+XCRwc8dWH0p2OZDe
oJ5UQgc8c11OzZ5GxkTFGrvaexGMrmq6vI4T+JbN34MPwMkx3QzOGfQ3smYPGxF77QFXrBC+AXMj
4qsL2F4Nr4busCG64vr4AbJAeOPHRBtFmLpBvFjvTwgjg+LDRmbmFU1OqeA3+Ajuf+Ifzb9MlaPw
ol2S6EYgkJ+xreqrpdJCSBRA+UJYgG0Sl2BEntWCfFwaVXqcGwHCyFFV8cL+kEelBpVPuB6APkEf
oVRF7htYZpWyzQRXxyXvIFiJBSed3ujco1ZOqhR/dGh4uusSzzpVmXu39hh4AGJ6U63d6k4d39r3
M7c8gvw5x2H2ay7cgpi2BgciIWJkw540W6sP5r8ej9lkC71QJR+xmglCSIq6d4NMuUrOE0APpw0r
YS6zZSaWhnIRdSm1Ee6OgeyfulfAujX2TuI9xqROw4F6KsSa8PW5/nXZlW/sK4h73JlhtF47odX/
F5g1iMtOjFu7q5Dz3GOm0UnzAxMbrapvkIyddBFzGNBZFQP2AGJIHyObiNGPgiK4u2vkd4zmM/2R
6rWwTKTsYsZWDaXBtYilB7lSHqyg7K0b/vYkOc7cniJzjV6kDQsWsmlTkK3A5CjFps8ejDAsmAl5
Tc0QQ/XmSY5LnTbtE2yZpjhRIq1HSlDCHRJpHBSVPuY6O9jQ/G66xpz6PeL2BqiQrLQzu9HJXvWO
kjRimmgKteDL43iSIAKsM92Vx7ZLQ9am5oPfU2+Bk3qpWzmjZmcaNHUjh+tsgI1HTzi3qs42EPr5
KAnLMIxSgs4DVgd9VF8GbnJ24RrRVLdXLWpII5pGN0/Sf4R4e765UXCpcZ3O3GWmih9axG6/Qz6b
if+OIsfCT2SsxjwmPaEbKw0jqwV5bSDeUR3d1yI106/Aa0oBh/crrm1CL8FoO6X/nrLS18FVdGK+
slM/tq8ItvxgwxYK3cCVDMy4crVDRDmFat8FGQNZyHFFvBklUG6CtKyWZ5Axx/BpJJNVi6q8AUTs
a2+s9gLFXltcHR0fiH64dIaghptud6ptK3EKxQ7RiGah6X3uJs665kI55AA2FECU5kbtZr67RPjI
QW/nMz9D44hKXYGjDpzbyHIMrnudLx42GdU/MSt5cpALD9LxiGeOW637uLtSbp75aXhYV3qnGWfG
fQnyxXgTQfcKUSMZbuwtGNHxxyG7CptliNblhgQyoOQTYYRmh/eViTFS5aQnm05p3QFzD8yPKuFO
qaCRwVT6f+uKQML6hqD5st9R9jJAlx0LxOjeLB0vO6C7QthLtp988ORPp7uoQGPaGszz6o3MiYMA
7PDPyTyJohD99ncIhpYu6ywcOcExQvfrAD6vMaieZ8kb1zinTvWVbdEmYa56bbyvV2wRcKsLE01D
yfOnZ/paFjOAFIlQU5p8PDvNEGV6VeIiZ4Swi2d8lHNuLoCIzaIx0hD3RbKli4Uk5l2kmlk66/0X
/mzLNqCG6vl0p/0Wv7oskbMmuXoEIIEmytA65vZiMX8tVmFpqjHGj29r6VVO+Dqw9XRK0uGmB9Hd
GSLtB+/s4RzyPIzadjQFCP8x1fc3VJE/CX9yM39QzAStMj1+ZlD+T5CV0+bwkbPNYlqQporrmZJy
w0jZt6fUSl/7BRl1GNdpzby22AlPW8DLBbxSb2RpCIaTLgDEeggDOETpYKSBqlvhqXIOanBF0bkQ
UP49oVlr0rQke64PkPswRhtdJWVuWl3XJ+rOBrfu+eqm9QYmnOLOeoK2lmsf56XwCaxM13/EwSPP
1kdNrCbnVxPtJ2aMDwv8aHvC3yhY83Wm44UedjhbIrR3lQpbTQ/nLtEYtyQtOKADbsC0oAHq/Eja
NNaAKpzJTw+z7Wc+3ALjRetnhMqUGaW9z/49cp7TACMvrGzhwMevVWPbGaQGWJj2zhnUPfTyt5kf
dfLv+c0uhtkmFLOBHAosJrL4ywQPAO2CWGUfOQaKiFVCkXE74dYnj4wEmtOwfELWRGrSuKCFIV7Q
V/y8O4et3nes5GkwpVUZl3DZ04MpUxLVxPHbnS5sx/jCLjqbIRXktUCUqQi0qomeMyo82jYr3gpH
srtYDsYwVu6uds/kiXz8olq+K3z0gdF2uAFWQvnQk9xxz8Ed+hoF8mLadr6f7L84U4MSl2L3UuyY
QBSKy93o1ryadIEALS/cCddac6MJpp5EZhk2r5LmEW7Ze9/Cukf7qNyO64XewhNnrJbIUbUeAFBA
OKna3AQzTs2ULBeVwCO6mIiMqt9pJl2dVSGOc23M8HvGy4BVlmMbRsBLpXoEf13y8C0qIZT/7vzV
VXLnD89DTeyDqf0Y8zP9KjoVsM6DfYKX4HYdJ6VQ6osUXcUFNHONdtDXM2QiANVzOFi44a2dNTbm
yO3HKq4I9aBIQdp6YiqFcuMAj4mFfjRjpwWPJzyc97AM+S88GGGOEkPaYL4sWZQ9hGp78ROlqaDL
xx0yF/raJlfhUAtN652JHh3AkoJvfs1A+fpg7cb1N8g+nZsUYW6+WMV5VadTlkEsBdHQsSnk6S83
oLaQCQZlfv/xUEHr0eEGPbsJWAMovWaVMbzUa5pDSLh3uqI5HJzKSznwSYxsBJHLt0T9iZqnv4hM
ODC34cjt1+jbO9bPt9jNgJTEJfjETRCmwjylTAN71rtszY2NQc7rnQaVl8gq3VsWSZnUEqCel5mk
qqGfzgjDtjE5wUck03cc6UhIgoGP24YNSxMClnw1tFoT2mUx0c61pdXKSWU1yEbG1ImraXXEgyt/
hZhVVOlnliZ506I3B8nhutv7kujxT5MEgro1z0oHum3H1qiiuqdidoVLCn4zqcAe8EjPm63hSqjA
pXqBzV0Y+eS2GjnB4WgY6VLk13h1D1uyBITDYa83JYOSnhTXeljEJKyxhhn5x9z0iqLF9Q5ArtW0
VbeYpl/rWut6nKPE/H/390YfE+yjYaqUkN17dY+FK+BpCsGGeY2hQhTz2He1s/vUi+A9RlHpjpxI
h0mnJ3jFZBU66Kpo+GSjm8Sfpi4E+7oA+I6bgPxuz/yLG4FkIusEUX2QAu5w59NtxHU+jm2N1THL
mMK235+tfH5SKQW7MNiP1//eFimfXY8s35xyZpDBUbvhmE2VZdHVzrPHD2sIGNta+pX8LUzRXsPR
KYBqGeCe/CIL9aXGfYU7KsZbP/PXNp7b6qF1vFiz8x0mhg2CkMfmJhq8Jr0v4Liuc0+nt4I8SBRQ
tbLS07YJzTBZcZorftCAFnP8YiIYYIi7gPPZZ7LVIQr5MO50mHlP7dRyyrboJjlVUHBgMZ1uBG69
DqV0DOtq5TTIHVmb5OC00enEGjrGBFscdIttHN4pZaWud/xjc8Hjo3lI9/C6HJJ+eNXzvCLFBdo9
Vi7IiXIqeTlb0XXJPyMhXGoyF4d6kSky8KZHM7D+9PrwNpkvV5Af+O1BAajjNTeA+tumy2F2W6tI
ljBqYK6TYcQblPc3p0ujpxPXSgpgrmiSHRr06wpL/j54Y4JYJBMzoHsDuIlLImWT7JU6Ja77/ljs
XvQWgV3GsnCQuCuCUUm6eSiP/jpjdTwqS4AT8/V8kQZAaCCj2Wh8XNj3vNINOuzlPSSH6SMK2xzW
pnWM1wyKqTwhOMAa3BFSmeHpZoZMGGTUBl8/z49J8YW0KZA3zWrd93Xy5KPSa+Al/HXm3+IsEGji
5nej1/ParK2qtD580Ecnm5KnrAlgqweBtTI4I1M3DB5ioNvT4KyvQTqsqmUNsaUNBSrAJBER1JVF
B3dk3MPIev8edOZwlgsQfDJBT2G4zWNtpJwEloCvXuCi6bwOEO5MlmNS69Vyro09BRA6tQ+FtaV9
wkjRUY+HmF7JxNkmSc77nEuA7kLvXWbXGu383J7b2biwHbm9cYhYy0HnXjdRfcgFeMBRQSjIXaQY
hRFD122U4kY96TW6QyrW+uKOr0LRC02z4/uTb5PpUUgMlzZ3bssvnKMJMtSQORpVriu/a9f60ybb
0wOwEeLoEC1CVZXPDB1rj6m096iWFfLTMNBq/e8XOFXsnIuPCKHfIe4ctN8cRt8uud+C+xUr9Wqc
GH69dwimEmn6q9HFchUIy6JW0y60uEj9bcvxKl+FOTqkISH2V4v8olMgcBMRRTQbM//UCL2RhiZO
yQ1cSdFbd+KPLKeoWqL7vEcUl+p6d761tXiJM1yF1quHacw2I+RZHLvAWuw2FvjqcNgbEv6wnzFC
UbFdLAyC9H1Xl348TSHc3bameDd1CTAD/r4YoA5TAmmUVDo/cbI2jIjlayCeTwahPSx1pR4Vejew
Bf7iUiEWLwxs4b5Sfd8DtuN/h1FebDV/Aq9v8P1P86qP02TbyIvQsHjCv00I1KlGFae7TXuhi1gs
17zCK7eXAFeL1PnPr875iYz0NpsVWSubpluyLi3qo1SZHl+imX05zcf/Wdjk5IsPqgsoGBFf1WYt
GEgPRLsft4Abuq1UjYXCn11Fk1KquCDH3ow9GyNVwRFdD0FOq1iQlLxZ/fMBP/fyFnbIb6u3PgxX
nDmfP6ZoMLqte32xS7w+bnH7+rjiXajSAdpMxrBnQIN03ut96Dk1XRtr06cyGeu3gwng3G5Mw/EN
/ehlHK1USOT/Odtb/AdKvkcjSGiW4ISYX3cH6pPPGgMwviaRM26NyFyrnLDIsA1pwVsBUVIxLKkY
vG3Vm3luICvJMomS3ZcsgoZ5DcXLrc0Mdx49QtHMelnDkJuQBTdlBLwz5kIPkP08hFQkD8sb9fqg
cm9C+PxciLHnIy7tMkf866qNNkIIm3xpXMTAs4DYyeWzn4rMPXridhteAJZd0G3OhquGiwIebvkL
Xgwf0Nqsj7w619La+A3mZR6HlRGpuToW74BEfC4cL1H8cnidOamdL1B/pwINbWvx2qksBPteBTav
23XT9KgOk+ClbUxfwXb7UjUFmaUfZZMXRLJ+kiZBKnBh5DXeEqS1eteFWTuhfc5C3FMLFgM3j7cq
MR6A+f8UOfkQS829W2sYTgpfFXZVxml/W4JU3o+peaQ++r5fwM83VJm1sCsnzGKx94hMtTiX+yp8
3BhMZPOYQTgpwEBItAXG80bhQuIlHdE6rDZJYw0PJ7wnH+E0fyvm8fR/LsTdbSsOrBYlU2ka+dnE
muxXBhiwf0z1jCQ+ZgphA3tK/GdB/w4SIo48DoZcke/uMF4ciHW6+HJ8xz1m/3z26wEOuvUhp+j9
YAbkibbhC3zzKYdRo+EcuoJ2/6DLHkDtKR7rUH/50X07q3iNM7oVlCuqYttqgH1iPkdOw1gry07v
EJmjjmFBtbK/hQa3IOG/bvSl0pTgoi+ZCbJc1YhSQCBth7kqhQWRl6D7Ufx2xz7ztfH5OqR09CKo
kf6DzYv/9zp1LQGR8LjLwd5Q5qjMkmI9dr7GeRNtGZEMGvxsrbS/wsKaCD3jPuTaginX4aEvKihB
XVElwakTsejXvhaQJ/huzP2LWFpmOcv3EuYa5eLExmO6OBxUvlXdUAc35uBLkiUnN3nZxLEQvop4
e10Zk1wBILfUhy0L5er1hj+aIra6ALNbDSksxLso9maxaoMeyaXdLTiiZj67jtqfafrE8kkOE/aK
fBydW0GxztNNBUYfs9Nbyrr5FtaX6ak20f93WIql1F5GMqgLKBUkJOSGBXDSRUxHuKjuISUG3R+L
3FrBZUqU35qg/CdRMpngDOKHmguqTkJu9Tvk2513pR8G/H3omslyC0qOVKedjDt8s9f/zLjATs7b
ZuUPdjBGXIVmZHdNTaZ0etfV5XmjYnHM5dyFpmpKSoqHlXGHgEFZPGnFHJ7RqcnqmegbZSGq7fZX
oJkP42NRt6JESO34SqTffxNEmVWrP3wf6G/PfLSMU57t3lBRTqBfh5PCUE5YJ0awk8TfMw02xONX
iArkXNAIta6IkZbW2xwGBYzHpDDVlAVYjEQG6BdJUidKzaw/z7k3O6ipmbZqZXFaXwYZJWs3SPHs
STuru4h+lMHqN5nBfD2rh7XZ9cS/BkctqPMuS1T7ij/T65SIx5u9RM/Tr65NWToR4TXfRRXLpvXF
AqbZAx0U23HKwRsftY3aGwf+edg370ssMyemv8u8NX+dPK5iPDkNQEoMF+s4xXk+drsYHJLQ4SU8
6+2qZNcbXkBpG/5IEiogWHlm1PtFY+NTegnH2CqhJbaCBeKGJdzGNcRdrRmMUZLWdgIfLD9St7z9
vAOmNYwbh6EbhoLX2RzGHkUqkQO1LD1TPif0ADwcu2xiulnJ4HOk1WJ7Ffw0oPg5UguaJhLoYSvG
EofObnOB7vayc4hXUkOp3L6Goqc8RmINYFTZ1tmbAjzA42Hr7QDFiVnRfj75eKAqDExEKLBPCQf3
Jrsbw/msa6hYkBEUe0WII0xUUqJtAYS3raZuYWoj2gQ0OTvWJ+CcrzhxF49Chmm88IZiHW85a6qq
GF5qTKuYnWBJ7ek7Gmr0Sg4dbOhrs28PyX/4Bg3qiAlBTzAvWu9K0k55cU4ZU9kBG/pqo8xbISDH
4bqnbphG3pwlyU3U2rK8gbLdj/yBFAFjHhKKB8jp6yo9ycW6GWmIDKJXy5J6TYE2NlHIatf1G7Uh
h75IKrqPYfj5Xb0LPpL6pidOsjuFcXvAiWNExwLmy0ztm/rbZUz2m4PbQ5FoJArNAk+P1VUUNrFf
bmRuGXD2/ofj7sR3PXoaRiQga1uL6RUpr+KfZavhvHxfA1SzdGi8zVdCMDT5ozwRVc9flMZQcKxj
hcGLlBGADLGnd6s5aaSusB75PWJ7NQHmxDei34L0bbXmysdfrKWElb32tW3yw0wh7kA8vBq/Nn3h
cUpdy5oBr0IiM0hcEG1bgmfeNStVKxfA0yaSUryvoT/xgMGZhsqYaWOBFP7HxNFgZ2mZPaar9RZ3
ZaLMcCbXoV+sBrRs68S3xF3emAMTPsq/u8uWtEhCRRRqXKk0hNxhuBWOn5+Wv8nzH1wL0FVN6o4i
qE2Fdikr75Z0dM3I/KJJq3Wf9iepkE/cfkIGcxOc97QLNTQRY5VGzHrEL3rcCQ6Lxr4RV+Es3TBc
IjCOUzC3Ysrq/qDVNDwMi135GsKmdeN1ph9xm76a4B6RWvWTG3iiLNMSOV/+N8DzlJEuYrT9kVfG
TxLVAKwtcKR1QPVNQC1jSygH/GB9ehFx3Dft9iayc9AI2YgXZkTyRsVLANqEfaDJWKn96C2VHP+e
eA3YdT4gD0S3h4ZNj1Tbn9MnlupEpA31Q8MvOXQJLuU4XCGeC0Q11G+XRGLOpGGD1OEN7b5euip+
yTOMkZP2j7q+qh9m4ahHXaH1JgYZlLvmeX9gAG5C+nYDIlFX1YM2ILG0E/W5P+9wgLsKZG9FDjky
f6H9JGD6jHRBPHfi1PvEotcNEtqCo8Bq0Q3+5E+9WcS1/YLySPUYnEaR4+1GDoFXYura55XXUC1g
dLlQlXy1DuKf77y+ZJ+SDRHrX6jg+oJyDTokXGAqeHs1BR9u4wT/fzWNmh7ZDJaIaZg64S78Y9Sl
2NajbCV4GBQ8YLKLqJ+OOtypx6BqB4SVWaj5X1bfSDtmv8L7miUD/6XjMfZWWN4PHUJUfYkTveVd
gmOxp9SGeGQfr+ZbSZjGzdaUOMgdwmUL5RQoT5vjV/dYO5buxyD6NrHgS+XtW0HS8lEbV0706LKT
ONMReCmorADTIl/7GP3mDAWsUWrlTkCvNT4YeuKM2qYMRBekykrXs933+k7x+7cpR4bYR8sLN7S6
BrcN26gBTVW4zKD+dvAO/MBG8KYV168G8ilNk8R80HhlWsGsjxupGArHfc8jIvZr9NqYnxolILWE
GP78j5Z3Zt7h7POF9+Mu5lEc1hWPr91RMhh57MCRkBHEszdoVpsYjZtdN2ApaVUdK+U594wBSHh+
jNVe100hVuqa0VnqRf/R3Pyzw8EYQYRzcz9qH3IN0SZx7kfx+mKs4gHApqodU9uIh3IYmQ7MtBRQ
9zwKBXhdUkMQhxHV3dnunEc0lzSVR698NPDe8IByhVt/aA7lHfw9alf++Uo9Vl09Zph5mqC7skWG
FxoIlIMJonseeB+sEgZ4GVTHeusEQRGJCs2lfXdBkGD7KUX99vsNXyDl5HVFAvtvt77FIj314Q5U
RCMMamSbLo0enuigflFxn/M1BcSx12WhyXRFEbxgi0AxXE847ltWK4/0PpHJdj/mpQ6qPahfzbXx
zsMxyPCQ8vQ8SKZMuFq3bAnRvRl3pPyYpuZWF3yObJjqah+yQHlOfa00GNyCZ7dcns0WjpTzGXn9
CwlKfDMLJQBhY/LArR7WzfqAR6LuIbaTgPVSQ5IkQxfGcNqRQvXln/Bi6/Bi+hyCB6YcU0VJRInw
wZkplneoTFAXLyIdhj3hEFqEpha7LlMiuDSXdJNtET7SUXv+CHNSQu6wF0+HWxRj4pGIOLHsf2Qp
sYpEe/weeRkzDhDEEX6eS4udllZIVQxqL0+rbc60w9W9+XzpFQsIEEac+vuOQpzw+tP4lRJWcFn7
AGo97hrImlYkq2NmAjUikCXM7Ui0gIQ2CqWgzDZ5EiLlSm8y/NV3WtIvl1DZ6Ggir86nrcjd06N4
U0DXmYTEE4UijZy4kZCC5xil+4e95t86mcY1gNLl8H2S8RvOK3bg9Zk7f7btV2f34k0bmGtIwISh
vc+evRR0aNbqCbsQQIgZ9bJ/r9oKQCrQ/eNrzcJEMmF2rTMcJE+rMbNSCnJdUnxWe3tLVjzHfUiv
oI0iOeYCAJu6Ka3w+vSuXR3oAtm1DQxLTOzL7XMuDWPX1GcLow2u0mlIpqtXjVCncGY5K62KJwS6
/06C+CqUYIV37gSSCdlMyET8U+UhgClDc2Z+DzqJf1POFDPDqEBe/1N+4JGpWRzXgm7mE6gKABfB
EO3mWnkhSPuz0laZUZy6fb7L2ZuUkfQ2NfCSboaBKkHslcEQOvdivfVKZwpPKYnXuxLSC63jGGx4
eV+ursqdMhasSM2qdj9V1C2hgMUMhc2oEowQNUItpyjADZLGYZUIR/tU0Grlko2HW6Crk5IkQEIj
MHjh3eNZpK7x47Qvca+yFoU8hJWRcStM2fYqsPQE0LxYL7rU2iZOCaNS+nHv7ErPG3sk3yN0pEtE
wMyZbdl5M6oxIXh3Z63ZFFAVgUfBS7hMDCdN+nXTfQsLj85XxW/H5wGSLPe4mCF8ri+O5v5EdxdH
j56+eSTnTiV4ZbDaJrRsZq6DUbrXcY3x2W5eBPICYMaO0Fcaws4EF/04pKOFMrXJrl+gewPd1evy
Y4k5sMNM3YYW/Izs7cGgfxRXyFmJUzGd3BP+q7EmfIfeVJ2lGqnXpIjcUvR5LFpwGahn7ekUmmDV
ibCCNiG+1X0us93rQRpgX65/Kp4hO2Fhtl4dws9rFH1lPj02UNEcrUoZVP0pExIhBZN5p1kbnSYP
2Dpd1og6lc13V+jhlVV/mrgrvOPOT7h2PVbJyyxCHZx3BigP4WukPRXtbRaPKRYi77sgb4eW/+vU
5j/7xLX0F2YVphKfebo0v/sFm9yC1KxAYIbzE9miKJBADt77LkAHQRZQmk7ZOJ53u0dQ+kzV9m2r
ig5yBJVSE+kywirxf++8dncPSJJUbg+YXChiYbn/JSoar/HGJbJe0yLCrVrKO0vP0a0CGPO+lzI6
GtTunRDmHTao2rcBcLx436kIPI0vBi7ozc8FnbjPqEgOtQhLVX1ZS0T4FOoC/m3DGmsXClsChawy
nzOq+fHSgKLFi1LfRsmFeyHQqtCUhGqUsINZKmco2ZV4vh+ajPshSSbd65WBYvbw1WG2Nr/zJL7L
2Gg4sk/h44DxvFwu7hBR9fST+NF7GlmIgDx5aVGGeyvQoWA/NSp86lc2rDe4N0WU6PZbyBlNUiVB
rHCzKt5sIJ/S2rpv86my/KV9Urq5IBeXU6TinECozdx+/qAOW0VrEj3iveD9ukP3rRH8m5wUkf1J
qW0VF0fqTTbZKA7Zr3iqbh1U5MNAfkVBDCJjQFO84zW2jgmUMsd8n02obWRD3jcLA9TpwkLxyLgc
/qrQA50IFBRfV2q38zG7qZTVKg4LHUd5xUOkzXGzNsl5mmLp9YcOjrLyh2DgQ3YL06gCy5P6wofn
lHDgxBO+BAJOnOu98mk0N993o8jDcr6suIYeQYH50vx+HKKN7vcjwjkuK69GmeMdgrG+QxaIavjT
LBQ+RfpjAjSeTbB8zU77ps4rbb4NBkJu7olxw7s6n20BvHwzC8qqtpc+SQKvZe0/SX0gx02sEyND
MwMUQcRm7CEMoOlKX9Wmzpa5+X7km3EhDR6/rZW1MFi+/BaMRwZJJLBoAokm0bKYMOU77XIP0ESQ
1U6v0nDCZ+q7H73t3lmmLcZSiUuZ8Pt9XcEZepArMhdU6LspIVNDF0PU8WP7JOPZhu80ovop3xFl
u66BHU686GPDyUce3GmaEWfWsZqYELPbSqlZtUSI6wOtkdcAlL7WlStSnKLGszNSIUjHlhrp+Dia
IyOskUqAm0N3sR/rGGd/goYjj+PAT2vUjxz6yZFHNTBbId4V2u369SiXeojUvxR/1K1CxR2Z1h21
s8IxBVxjGDcCwyqxJGH8rYyXUQRvOdnPJ0rJ9/4vYuWizk2cYzcAjPDrMr1AVG37C+1azqFbvrM7
s8Ik70Pxn5QcZnpcHdJRIZi7duo+LytAOGJlYRUbNE1s1Pq35L/PBrofsoN/c4fvsRAxzKdRxjRA
ZDPK23fyfD3C5uBHAQaXsHR2IRYoRNcf/lkBM0iGUUk6YbSMLZJ2EqO+rsS8VMcXagxs1uqC1Hek
sGwQaGKvwQcW2DiSWndCKX+hy8j6W0TugHB01tWpt+ulL+SGyiwSY4YZfEGz0v8h/MIXLCdBpmvW
UXwWqrJsnn7qWPyRUt5XQ8MTl5OuAxwLMwnXid8TOrxcPzQwc/b8sChkIMvfxYArrDlT0T6VIfk4
s2Aj7bkGttf8Z4Ee5917OvVmbtYX6M7xE4aJFqo3MBc8zNWR4ojtxkKrOcvzH0xMkj9OG+4TLdAN
QvT09vhOjmst9apjRmuaA2HMV3g4QA+2oK2vPEg04cDATEd3RPPd7pYm57abXqK1BGyERR18arjv
IY0PDqk9/NcxTGI9KJNRuDgc9WVCstj+HhHOHd1rPjrQHjklqVxtO4mtyevnti6bgQDqvOmP0o+O
82NW8opm88LJ0KzKcSC8Zn2f3bboFsWp43JLmIx+TfvWWMbR/PHvpTFWNyH/T8QgEgjq5Z8ONtic
gyUp980j5Bt9a8h2A4zYRTDAoqBt5AJM19TQe3hekBspFhOCH8YTsCJqbHIHoyvOfB9cimTMvkZo
qOLczxZLqa+wgq2FZrdys86t59dR/0cllHMrbLINkIWbdtOOiuA3OfZLcnWtzVGX0W0B21cwZdAb
O66cQYnerU2O4sQC+CbzCU9hAZi5W0Ic5htPWcBUCN/yb3wxSmMof+UIfIEyV3pIQVVco7BtgJxR
IH01X4+fErxNhJDVbIxWYdNp4V5l6XHjLIHfjyxRQQ0Z0HO0UKsfhLQPJTQj9AUABOXb72VyWl8O
bCxktMRERjKyLpVus0Q1mlV9/9Ro+O+DMbVSMsTFjp1K7vx/SKZRUfDJaHc8FMSxbPBB1nMij8pv
jwK4kDN2DkVdk1HefF1c5PC0KqkkZVpaOCXw0Ik9oxXRzuFhzAc4488SF2wxP1Yd5bYz8nNqkylV
UOcf5ZeeV5vV2a1Fca/RZLZC94UC3Dj1ibUgEIbcHqYQbKvLoKqEG+EKv9Iq91YZVRHXIPPPrTCF
t0jJXFyzlFBthT0Lrtf0OJS3FHmR/lu8JY51g/+KJyeNevyBR7B9XA7TConbc+/c5E1DxEkGR5gz
9+O/sEog3AXcgiBZD35SAXjz2Pv/Zbh95Qy/7neN8qQYIWsZb2lKBK9ELgVUw4W5sra87EVwk8ph
sADvEAo8tm/+kJNLIXXrNcXUgzFdzZaj4xY1QsbAm9NUWX20tatNIh0x400+yxgjoOKYelESYyoI
xUWI2uC7yTafTw6kTPbjeDg+DDBm5b7bvRfI6fI7i2DuYj23dfYeYucijiQZANwQCFF0qe2Xpcc0
kKQHqTZ6bEO+DSIHCUT3mBbZdpnG1qz3fLEAdvtTXJxUCaV6jVePvLn6qEsUP2/AqWil5uXBfHzK
qyYNvRZNBexJVa66w/G6EXX552dgkdx2IVu7VTRAiXh3/BQcQ2qzTqoNSkugZz6KSK4xX4NhlyVU
MM/OYfo+ZpzjvP/miv8nR5rl0L5us31N2zqMmp6o+CtfOqyaYjN6bW80d2ytyLtPnNyf7KnxOZsc
7qsRjpiNnWs/Szg488RrD6IFl7YYqoGl3uU7cUxTJV8t+/5gV4OV/GiHKgBLYsK09LDdUu+fCP4u
bQB2LJuGB4MK6wqaF63lqy2bp7bHSnGCpjMg9IbyR2mLndgVXDMKn61I4jm0fxmZZd59hn7YHhiv
1gH5C6zupEHHFy6krs4FunOItpdkkC+sOj99bFFeUdyugUkZmBXVflyzxN5xaZQAZB114oDYkCb8
QxDsdwyCwLs/wHtzgmarxOIxj+BzTy+jN6MNtf8Yc3U4wVKTNfHzOdbNn2ONyJu/3MLrtEhk1h1N
Dj0ozxjXST1/G7YPZ6oTtvY/kMoNBMePeHklCGkwlXctFsNCN+w8Lt+Ox+igqdV/w8inMz8nLxT0
o7xsVIY+xcFBLJPno8D/TGO4dnkzjZc8evELh9Z6d6HXzWrq09a6uvnxRKxjGn1YBSiXtaECdDlB
FsTeHQFmCt/K0yBgsBMaJK0RbdhaqqUSjgv4/YVLLQjtxLAJm3/nJ3YRIwy2P7rxkN6YFTzjuAYp
KYxgRFJ6AH/8PtNXIWisN4bLqcYr93n70GuglGXR3xMirp9qRpWWe6alTEzDTZntXtbUyayXaaqj
es+DC4i6FReJnL9fnVrUn+R2hbDpyuSEhWTnqiVBe6TfU5vNMS+g0DxRxp11A7+R8Znv2WPt521z
NX3QE0tVLAZUvjhYx9IemC0l3Y4I1gkx3eZQn6MbCtG/umFrpYF283ovfEMIuFeJAQuAhxHsdMvW
fLb2ZpLpQK/83fgGdcaVU6hwCQdwgPCIWu2z/6jVopqQG6kw2da8S0MXpZ93QbSwJUw+FAzgVjWa
0SiDa3XTTogW62ixQrtd1Y6Rv5ErYOHrU8JTvyEosqsqMWIl+dqahwbFkATPhTC4Ml5SBQka2XQI
SYRqS1kRefGZGPkYLCBu4sQ4Z78kj5lQ+SwKYHQke/jESih8mlkeNVpLdO9wr7ckdVuPNZDNsuMV
/+n0Cp7OZ+lN9r9oWuGU1uBf7+A3HYkJmkxKoi8b+YQWoOikMkpRb+y5zuE6/q0BTNmw6G8Gi9W6
WIoLxNrIwKOTEb+q7MNGnUFd+BpMbpico6ESptIFx/weVfK7hQICGK9YGvmcfVtPn1sr7IfyxGRK
5uhrrWjDdhu538ysOQV09Nk9ROeL4lUaMdORbj+4Fw/FbtLBCpu/BQTQQ/Fzpmr3taXXSFcBIXEF
qx41lYkLmRzr1GaOEeS7no2XR3OvGvEx7HtCwk9LQMQnE7WHRUZ7yohvO4NcsFnBPu8DZJtJT9fl
QDhvux6/Hqasnew4OIeXMM+19LZSbQXoe8MjmPsUkB095kJp4UTziI0QfelpH341SXMisropfR7A
8348mmKUvu/TJGQBkPcRBVTm0HfpCLX2ANpkOAzc0xfaRCAXHoCqIYEMyq9jlL7XnLoSjAYR6NCJ
drFx9jeW6XvaEVEiFDNTBIY6Hgd67gmPS//AwRK4fXNYVEfF1axcgpiMuSE9Z791NESpawcz/7Y6
cGpVO0v5gDWd1zylpTBXeU7r/dHE5I5nZZPbgX2sbXSNxD0DL9VAVePVO6x4YPZVpzWQ0FBDJeT/
Nc2rtaHGZHjXH8y5XmtsLAK9AHdSVIxaNzecGbJfx22mN9RkMNdBFL6SPgXKd9kxwrI9oCnGV+JO
hhBfjJsanbC5pviZNwuXKcCLr8oe2nQAaMrur9+P6C52H47LBv9+JUESOVVmr902jKe2EJNx/dEQ
RYwmfEbF6wpGEVbgPr14ODdY83hWYMPcEfOn9Wm1ikGpMQhCzT5odQYbnETlfSRJ2kBKgF7odWsm
qFWa86xUIsaNedpLk7/UNVb4wKNn7ObvVhMlbFgPg4dDZlunfEJhKsKyBbjVNYX/RFZ/KcqY8VM3
7h0/a4BXSpZddrYGuNeUTWhjeC+EcigDwfR6RhiUh93nEa9w0E3UAxwOCYG+p/NAZ8V4Z6bXpXUa
EdN9ZgHi5OD/AD4uK5EdMlaeg9Cs+4+UhJEonC15FGK5V6qPY2s41g/kVjbp6jpSvaWsH1cDi0NB
MwzZ7j36JQGQmpmA5imPYA4VglEYfNpBLM0QzcPMFHmzvalaDWe1IkwRK8BU59cvrH2dR7CqcAeq
5mpgs3exsD6SxoU558atUIJ6JPE1y1WEi/ejaR4eXmo+8mbrKAqti3uoKvcUwKKfMoAKQ4mNE4S6
veRUS6c+qHwjK701RmZs+FlXioHCCnloDi9UttLwrapb3hvMnCxCN8ip9TN31JCHo7RWSBbxoEHY
JymPjlfbH2wLrKi0Iq44az3w+/E/TGGNGw0ZY1mYrdznlm6EKzt7iNB5IbXgDiKLhowKNuctvB6d
4ZTNWHQSfI7wzovQhevrKBQgzVzXHdemoN1lXXZeGnq5fObjRAxOHC6m72gU3c5KSt87k4Gm0wnJ
jiaLCYVrlNiruvaCtyhmp/BuKtt1mhWlvW5YlAj1FuDgHzkQwhBjS57ffJyiwc+Zfgf8X+Evs1mT
E27UY6ol/ZZ9rR4DnbIe/boRLFTywsv3MDQckXeA9ox+z1+F02utuESJOGI8HBTydemQ55BrDA6P
Sqejk+ixD7BIlR5dObS3TLKwELulfqktO2gJxJU2yQEKiqzKoI+Qp0+NWH0iV/7//E8X7f0Eneeq
SmUfxMJeO+76VvKucwYwZHq3eXl469sTLRJ+1rZR0yg/kvBQ2aRGUtAtGNRAmZaWDypEcFEziKJU
DRa8Ne+OAzcRMcUNq/qsdomvciKD2vZ1gBL6suh9KQ5iM5ApGd0PUZf20TUFIWNCSYgJJytOFr7+
xfcq9tvCi2E/R8hE9KaFXeFksvjo1yfndSJLSA3kO8ivCGaDoMNbURp0Mrt8pYP5wTjEzzXTRs64
zOCjgeOPE0Sjb3omYoYzLC8bca/gHPUhKopBidxb7hJCZD5fhZH+JIxG5q9nk9tf8t1HIizdn8HR
NDricIdii4BXzfbF+G2nsxmby1l0W7hJWTG2VKumAnKZolHt8bB5SgVAdjWox4uNEKm+nTdD9YpY
bG+M4ORe9LMWn3W9Z6p4+CNegt8qRgTbbh/OkzZwIN6jqERZb6Aitq1BeGQOsLXsUkkE11UtsMWW
rhIswZotWiFVn+nHalO6508oJ9H65udXSS8DeoCOGsHlOPy+jwhDCuak2Wf3RyjK8Yq4FV0SUG6r
Bw/X7+ofpFGuyvqcuGyWNzHg2tlnuYnn1XJnJL4RixvkfxGKD8kINfP2g+t95rF3wqiToYir/YMl
OQdEJH3sdtIxh2oVlQhMUnsPG7ZrcTgO5YzGSI83CxyLa1qQFdQCqLLy2aNFTleFNck+8tQ2ELLp
CzxtCNwVSUGvhSn6W4+KzN+YEbktoSmBjvQthYXXp+EK+7HNnk7m2Fcaaj88k+DWC+4EJWb+bdv6
AHk8xvIpwuPZmS2m4oB1WNZBUjzAo3gEc2BVj28LjFwRV341ZJPMn46h5UJXMkoHRQfcaow6Y2QP
WIR6Z6eaf+S3rjQntUYFsiRLy8Gyjkm5KJxXLQzI/oQg+EST+6En8uGAZQyADFaWX1hJZjO51Weo
7fKglt3LTtQt9KL93nR5+G0gaSwGXtHyOX+LAauVQIuFJ51oSnhBSfZ77FJS4ewuu98gyDqqLDcO
ngPFQuKfzpbiT2hThQmjvayy8s7gQEaFShcasZwPjFRzeFfXIfL3q1BB5H1vxZ75jTFqlNt3HwEu
wPGTrUhzT6u1bgngmWYlPzCw0AxzSG9mf7uLGJ8MDopZtoAYeFkd6ykQqZ6w004xDQGeKwVuRrp2
5c0KA/JR85fdPPTCh/E7qEajSohhPXs7JjqJ/3iMxifg+RcYgHuceKdtUth4KP9PiGrHPF2EWPI8
W0eOZpD6VB+ZdZ596y6yucfcf7cya0bzdyytdhVdPCsnTaGWhf09kBCBOvgDeGOJHD115f3YlafY
4ka5FZO902Zrb9eCJTgBCaHpm8BOssoInKZqw8PxS8IP0SBJFEFozY2xDjCFOuvQOzyZ5yrZKMq5
oPlq2MYTnUh+2KIr6aLYb7jbG723PgXvF2uqnFTpHbcq1OPoW+b9z9bTSC2l4lHGHIu9+jLpHnTa
4/mD1XUHAXkIfg1RUsc8r/AQNHQURu61loG0vV6dCJhrL1Zqoyf8tJqf0mGBS9qFFA7n+6KWACfX
I3tcgXoFHNqRisxH2nRVTbf1t7um58ma9ykVT7zdzNmxn0epfBBt2BTpoXSsz6N9Y6d1ANaLTdb5
0EFntH3jhap+/VGkGIYDJ/Vyvy06qM0mT3ZcCHb2lNFxfCQipquNP4q6Fkml1Ik5ATeNUAczohGo
dlAEODq8AXdsKn0utirvd3vMn1s/SGtw0MksqmllWZoPh91032CGONQWkbeCw5VjHOStDcwoV37r
53PrLDGn5jaGY3IyN3UvQHepvzVanBCPqtf0wYSpgQHwRZhU2pzqaR1yTOzt0yWwTP4FeIlrsiwL
Y/IUVeEOEV+3Ul1p+NpcHMhXpgT4i7RWPz452TS0U1bDMg+p8WR6F3gvoFJ6AS1ybmOm1tTi7qkD
eiK78GlFVi5V2fqJ2cCEUvXNNGS59ejTtDZxBcMuw4F2Sg1e+yqIaiiWzH8ZBJBHIcMLs9tRFqfU
Crh95P6CoxlfGYe+QzHBXi02+A2TMVy4Q9W0qLsC6eTCvfON27it5iqw3hyrqhUWIRlWKLQVvoMw
k/cQ1+xV2HqMV09OeckJIZsuyfLMKtjzlKrlRxn/AsbdrpTvARMlVMlyc5Qs3iyPkmtA/b6pFMng
eeMJdf7FMfG/6J0Q0i738Lf1oDHIULRcPwbEOozfbe5I4TeRIxdWaODK3GTKSZj18TvtLkgDsUhb
y6joRKTQcmLRMnwOQvnjvp3k9FLJJN08gLmejPo0BooLNYQPl6LUkanNkCxtWGDJ+B5mUyAIZGoO
MCfFTo+R9W/yEyKvr1wphMt2SyxfoRtVZSpBhk5XFlbC7BrXvzePJuSM033aAUeQ5PQu0+ghCma6
l+5DP/CZQVmIKPs0VnCVxjmr8L+9MYHG2YXUc6mGuwmGFUWCD3nZ4zjuWyGZP7+SFWUlU6Q5oXLC
oYP03UUa04z4Mnu7B+C0i2adJYuSk4o7UaSvtHz8L7GINQxWPpGpYMr5MWwH/5S/xmDjz7ZwUC8l
S53i9/ARSmFYgZWoNu0NVMNeI8lBdMnHPcZuitRi3R2NDlqQHkOgnWP0ScQJswkFZKQd6iRoBNZI
0BQtLH3vhWzykRPfYJgPNxl5sfPN7VYZcoduud5/G/OowPImPGnVscouPu/GhfvVs4/9C5qBo6W6
c+vOcqSyxFNu7RCRYY9zdrcUueI+bTQjT7q7C/E8KJ9jApLPVXMV0Qbej/HS3nm4t5bUhhj60UsL
K+95O5teHY4Y3lOCmrAbMMDw5JsVW/WOXHUGP4egAxPCMwmVuhtaA0bV3A9Fyin73HVUgrlW7NTs
M9s2rjTGfXIUkQOlHBIUBzcw6NKSND3/M+buxJO6MB0lscUUcKWMce1+YZxB0FfH4yrkXrqaAb0O
KW5thGU0XXt0cBFg4Qu1pKtC+eCWk69ATgATcilyVanHHdlvzGKfMBwGE3rZ5ChKSPmBcXy01Qpf
EV5FNWmy3WY8w9p3EwTxJRvuJUPYjJKtFAz54a22ZO1Z48WTvNNFPtPdDXw41IjqtjF0+swbAsgd
smHL8UGHJlG+Yi0qmePNbBxS21cbFGs/X82nCWaXXjko/e78cVCB6gK2R2ofFYW0lvZkPU0uT1a6
LewoOtS2n8b/exEs5Wd6vBIkNF2ZH4zzduwRGPpjnGYa6/CNC10yhqTcxtBv6bhV9/X1BNMHdY9s
OgvMO4gXtzQAviOqkXV91b10sWZqpHFGec3nRZodPK8JdC9JczWT5m+jhWtnzb3GTAP1efxFE0nF
wEUvjupClPmE3IGsq/tIqIqTs/nuLSOcSiJrgjUMeEduIuq2bVig6cRnWjf/e/73R6O6fgqJ13er
EWcaPOzQg++XZapHBZ+DN/mYdQ22S32TEVBXQcnM1fKKPU+dq689SDx274vmnh+ZXr5M5SoWdc8Z
uJdvhX28hBcSJKSoKwOXPMD3rijcMGoJDBvLz7/OMz/Gzl/nc1HIWvB5BI2cAEz2VU3JU380sEzq
BahFVrPknARp0oxqz1vstiwqzJW6nfA/wyRH01aIEXE6DkEjn1fpCCnsVrp+K0kJybJk9PD6RZui
l9w8ZJfAiDXTQIGV37SooJn6u7uxT1nuBYk9xNihdplvr8yMzC1fp+kSD+npHr9UUoDVmtFFfJU5
WokNNzBi3y6P0kMHT0393wx+2ZN7hRxcdZfJzpTAyT5wQVP8fBV6aRcN6G5u2YB7diKqsOkUmD5B
7NeugWRBhLkCsxnLKYBe4EZKEU6wq+nZMUJoqYCUBqYM2IkP+/IlxeyrnPqGvV0ED+O/ZdAg0tUH
35f7cYH13NJYHN+JJfN/p/W1yXp78Do4CAY3zMzISR1XhCA1BX2AD50c0xsHWX9WIz1T319fayDK
jBaKB9wq2IRDLeWoXr9yfWoex1c2AkZq3t8sswniJAAODJg6lplgFvvqsR3ngbsax89ZZ/4HQ9Ce
gsK4oQ1zdlt0AJAJTCS6fQDGy6HapJBS6bG7HykpNXZFOIyTLrN5RIub7RZdubEXPgI12Iy46HtX
HsQkeVc2Iv9qVvRTWlm75B2X+WHUvpc8yoxuBJveFF75JbD1iLGVMqtaCakDQrO46I5YmqLyuME8
GjcG99u2i+QC43OTvqPTlPVBGDYlYWKPnQH4OwS9IADahu2SbX6mcqXh+W62RNyY4dd9jvKTn03H
R2o3Gihq57HLUqVCFjShhlz8BDFn73i+7srMyOvNvB2hsZYoVUFZTGCZ/M9YuQAcMGFhM3EeIo/3
KNeRF2Y15UX7SBaqDhWmM8Q5o4hYsD9LZQkzQ6i0QZEnYGJy1kMkFojMg/k/n0zMKfe48fcaAFUM
6XFwSaWNDm04UeGYyAOzBo2yFrHULNSPJO1SUL7zm10LVZDYYcezPsr2xn6F96tP56DKCM0CvE6z
Z0rre2+MSWjbQKPxRaj8/3TTVOghoS97T5oIc5zXDdrBfdMd/KrVrmiP/6k12l5lndlNP0MfikWy
pYo/cUflw9EWZ83bcDh9ymxrO2+gwh6Y558xy01zFL5k7LXxnJkUZ1XWv7HaWicsHZ2dcjK3X1/l
I4/QRhmOia/lfvAe+agwe4Ct3Zk+gof/bTxlxdt360HiFSkXz9e0y0Nj8s6BB9o0UF2eewpL/M3j
tgf0gO/76kNjzS0LMVhjNrfc06QZcecnPKMnopjZ3MPL5o6mOkmJelRHTsYoRWtUO/JblDc5S38H
m38lgG1vZvQ8SHKuLYS8FmR1GE6HrQ9OWLwl07F2Q7gYAbXv5zwNi7UHjt+HVvyP4Sbcq6jFNofv
NjwB+N+L4ZCJiycs/NmvMiB9FTaty+H6k9ypd7wzp5VoWrKRfd7KQoWuIlU63gNvZbBnugCgybbR
akKYcs/1KNMLQlC4CvylFf0r0vEKVDkvL6j11Bxmbk1MavZC9fLrSg6ARwbTRQ2gpjBmVM5B5FZp
vrB44NBRXPwCaIkSwkDN7TTjWE0yZyYI9GgQmJG6T/NWgPqaF4dakj95EEzaxWvlaAv2YlqzxXfZ
KtdxEh3LWLNbrhqCYOD7Q/6+4PWXSzYKBBUbUE+Sx45PKBMv//BtO2IQvuV2g9tOPiwA+QARUdZ9
zYP8LR0AgcDeH41EdiWLPm9/1TN8gYzRGAD4ikHuZ5yv7hFNYVkUPpjspTyI7KADCSmh5+cQ2oGq
Qwmm7PT7wAMxFax6IASAABT/+ADkmTgfuUuectQIN0/rUV4z7jPDIQbiY2WpjMu20kSu3rOunxJ1
A4Va3p+p+3HMMyTkwk9aASOhSu752iYQRp4IIJgK+N1zv5rFIWyZnM67XFevD9Ty9dgoqVyHhgr5
HvGogwDB6Dj1UqpCjXXztWTSC140Rz5X4Cw8hQMhO8wmsZEtXabpdBu+YyHT6bKonvbbTOw+3IbP
olp3pSae7p4jfFeaemw2jlatT64QqVci2vw/SttcQlVRNAX2Kzs2Te075W+ojupPBlHs4qFeWJ6T
YbYn+ixCEa3f9mq3bxSSkVBwVGMNCXzd/05I1uSNkch595SFGguAfffm7q5Jg2HsZGDtxpjPs7OO
AYnj4DwsMhslGPrb3eCVu5s8tT+hbCYNLSRwc8Mbrma2gtdw9kTQUFhMrwJR2fpQv288j1uDe2YD
N3Yi8bYewy5YQvC4jtYCI6WwON5q/mMDferazMVVVOMUqjGfw06dNe1cFIntMx4cLPYVrfGugyfE
vQRfEBcLTHlBIbpNhmEvMu2gth5+JXdNmzza9wSdH51es6/RqA1IqeOa6CyRz9oX2xNznj7FepUO
GevB6J6tTAIOPjSh8B1oV07bxmCHZoFBZjosho4d83i5mKKsR9o7CMl6OQoKkclLGiiWRoTCCKh7
DJ18E28PLsnFX/zlqegP4un8/uTXLeHFgZBCMaxBD5MI6X/oQrIpiy8536Jt0V5EzjUmYZsETYCU
fWGCCRmfoZqRKCTuaOTM2HtDCV5FLJVP0Q4ok1TlFmVFpF20E633mgI2CyjCLQqLJbDbUxd2mM7J
DROe7cEnkWzYiW7CKyXxRO9mjmhfRc5psb2Hr8RNTOXxke8zy/dF8rzP9aNPfW+L7UDjRkq03fSi
Qi/2//RdSBQPWlCVmYkgnDy/plnsWHn6IacU3SmANzlShL+aWIIuO7+6w0cVxOAcrwV01TsEhus4
yEbNxcvfeHHmkbl/4hjdiZoQXfrf5VZecHiyaSSjdHlRpmrO1rdz5MsNnBNCkWIg7sz2iSObFLs/
CfFI/RbN8mQ8gikMysdAcQDyQWKWIdwi8+x/+BNMKu4elSkGul4izZzhZUhB77U6K4iy8bKMEvn9
LofECEvAkbOkA7DzWAjkdI8gV76k/TDQI7LvvGVUQL+nqcPKP/eTpRKskT92MJluWc2CyES5c0z8
7VymIWOj/A9h7Je0DoOkfTVaVEN4cIrOAuwDj14yA5XVRVYVW/WvaBgEWQ6gBledxjOMn2TdvRPV
BqfEQgetb657gmV2Xs+Ftt8dj1+MoDuHxAVjcmcfSSuHtfscmjhFD91+nJM2MjxofOxngqu8abpj
cR8FqHHn4Ubg11P2QsuPYC3wJ8hwBC7HHhWHpCgzE+JPMNJu/R+A26/dDKVYPvi/zugHgVYY3Zjc
ZTrA/iEx1//6gAt3T95d30fbZajvy549o6CjVLjfrqpowbyC0d3f7rJNHklDPWKvdC5NsnQZtNtm
wm7x/cdmIXDffEsbb4ivLuik0bj7TSH1Qv9ROy4mKH8yP9+LmQWWdjxYrLNrqoC892LN50JCDLG8
EMsK/XDDxWApuP3g7Aat1MTdsFTS9ptKjocy8Nx4vQ6bobyXAvC1AV38JGL6WH3/ml1A7p09slN1
e/yGQhJxgGa/8TpCYtX3oXvYTCjmbIrQ8Tx2Zue8/LsI72VE2QErU0rKquugP1DSvhr8/fTJ34bp
SzLaZ0Es8Uy/PqKc9JfVsJk8FDBsUcf4h8YZ4EM2oYqCfzySL6W1HYjsRQp3FaPXK8i11N7teiVe
4HRaEhddgXrzIEAlV4OHB3Gaa77sJhUD3etQJAdVmBqcBhM5MRlLXifahe3XlZCWfVXyGfK0MYpq
R0O7Raj/vD+6rZGKhusuxAv7TFsJjHxFihTriDyP4shNxjYrHyBzzSP8TQr4uYpQjPvRcjDHBQbH
iWfRMoqQd+5jPhiNTt1zhGFMEBH+JXLvZfvzNRa/vWnWvJwNLh4Ow5A8L2DED85Ls8Xmf35pYehf
SoVnbx+5tlJo8SnG1ujyjzmGZ7caZf8evqyIlzT7XWRtOHNvixD8oIRhzGta+eDRgKhVGS7rrhH9
7Jc7WVj1o03cjmiGkcCIYAfOYGDlDWYIRZGgKdBC+MI6J4rMgm1Y65abfpOz2LH2YLrcrafm9G2P
5DLni2aO1yHu/UrmVFXK0eEOl7WnRwP5orBsTLrsUBd6Lq5yUjwCDaqEDtUybmtegGGpS7IhFSry
GAAQEDDIOAWOBS7unclPLqCrq7Ja72jhfGuEkltxAenVBlHVHN/0+lwqEz6bZYfgYUUt5JuSy89y
aAyIqbrXZcZOeJSjio8/YI/208QvdVw1j16zigUSuWtuntiQEP7yisQcGDF8bzNoKR9oUMBOMdsG
mFMOlEg3OA+UNkGdLK67prN3xjsA98Fga7u0A1v8jURPztFK3ZLnEgk2KmEU0m8ml/+nXsQTouVt
p4Cx+xzJGbvW62UgZqCKZcEPNFYOZf0pp5ZzBV22lYUkgCtWtRdSdNOj1x/Ic+ApedXJaZfoWqqB
/Uii90n69KUq0Y8JpRp8J5zfH5Ur11FAWcZdigOCR9sYZjyXlCnaQ45gIfClgyv3VilDdVbrSzpb
gI8xczyhX+Q6L5KHdv+FxIl/y45qFBKqSKfZt7x/SLS2qX8FsNHobWzixVASPRts4LRUqQU1+VKU
z2wd+xRto6cEneGUO4dAHRGoWAJvRR3CkxV+ozjBt/eMiu0fEft2AtyX/NExHeERDLd7uIKL+axq
u6LKAwccspM1O9qrKwrLAAFJ0CFmROEjkL/T1IBAdP7GhV0XmFmHrTVpYylOTW4v+4X2d+9cng/M
vYdbA0sMh7SnvBqsuAQzLDoAFh+snE/ktCNzsHQE+ZnOkBa8n3FE6W9obHuvPGlyyCov55adYIF6
y81jYMJjv4CXn8f/zL+kpxc6PcmT0dlcn+opxLwzViZwSBk5c+y0+UWGnt+Nquf0YUTASXA6SDZ8
EqI+j3dVKhZgX98GOI8Wn0CosL8pmgg6g8sDh6nm3aUOGdGzCkjSSrMHW1wEuxO0Dbb2CDFpm83o
sFOq78U5Y944IIFrCXI8uUXf9xonYXwJetZM/Plmacbxc9eyr+VZlIHFSV/JXnOXPp0aVWGqlBsC
SaJFym7NvkzY2RpW9hpzxEGUHfAPr9NnQB6fiAg679tWN3lpumZ5iM39shwipiqm2yoHwHstI2nD
/+4PcXvbroQx+ReMSrKFYyrQSJ4eRnnW+cgMOu5iv+EY6NI+WUz0bHQXWBFL/c7Yi/6Tdtf46LPK
GvUWlg0Y1sThMHf7Mfex2yz1YNB43R7oSOu0m3yd3isaF6k4Qs6e27JtIK46ZDi/YSBVfHUnmMw/
OwYSfBTXT5g7y9XLo8aR6OOMiST6NCKBCmW6bUH4CsIRnuKu23g6gHaW/a9Mn1Eb+X4PkPeasAWn
fal9WzDY37S/CVkeUYLB/e/AQTGgMdT2V1Z3oAvEbN9P2p4glXPWH7ZMyXgE2umVGqhulchg/ixO
wIpQ1ezMW0cROkHxCPZEoVrluDIqB0ivkFc5QQHrB56Pom9PgmFDth3H6UCa6jQlNSxkwamCBSb7
0kcVoQG44BxW66Q9D8zkZuCKRZ3tn3nnxBRkweNbZn5iJ+0Mr2M3c3WTHCo9c3rbzIigQxTycGJk
8n/zcLlG3RXVYIORD2CDZC9/sEpdg7/WR0eVkB40Rs0417tOv96Zj7jP3FylQ60L+2DqCcYwL+mZ
emj+/EWNsobMphBV3W3G91vPovhGaWQCZxDM8ijxbPbcPd/4ja9zz70W+rCQk9tWNCSA9upKBzwx
tS/Wr9fw2qtte7dwTaeW50jx4B8nsJld/rN+M86pt8y4c6B4njM8b94vVGi1FWtnSzEw7kLvP0hr
c6LSdlAU4tOAHszUGhaKnYErdjlpjWyFiD9bX9TIECIo9bHhE3lw+HLbst7XRFGcU7ES86ZfH7sr
HbaqAbVgGCZ6oY7qgc7MW8m2gctHt2jB9H0Jp8bfaCH97DMi1h0LSMQriNUHd5ybMrjflVt0oMyw
dvFxxDFzXFkCnIzFR0zm/GpT8/K59rCAfkKxyfRQeCRuWhetb6PKicHpmk2wHK1PyG7q1ycPAQNd
aJhxhtqg2SpNbTu/mACnetxOZWbOUxDb6LZTE9KRVp8qDOVzKIrgiozwloHBT0lNC+mgVbnIq+PW
aa97BnPwUR2ukl+5MejAywDMD1BhgBV/dPpSKceYt0j3MjGBl3os5i+7+LG1NVIdSVt8nKF46H3M
COZTXQTPrMwUi2IQimmckJEEdh6pWAyUELPEH4xBlZwOFSGLWo7ei/HAjP+CVc8OGpPlG0+m8CHD
G6iQ9cRgUCKJ19CM0tg+GeusJ3sFR7HuIqxI2zIvN2uJ5ZTP6ehRGhgsOZXPmj0FRIWXSOsnp1Tw
MZ4ajM6exuhmFJBCOo902on8cthYzsRlGL2R/UI3Ry9n4efCOZa5wseehb5mzD6+J1tBSl20BvG1
EsA/sgfwRlbB37Eks1sfwIGaHKO0bmu+DZk5TMixvUrrNK1DJNparjyG0MQ16Ujq9KnDDVUUgXao
62KkDyMUjjDzsYlJ8xxaudk6ccn2m8/0cvSZxONjbsB2sqvVyqVFS4k27fzfJ/Co+8eoXwFcPb+i
edVlY5awznnGJb/Ek+5FWoDJNZpHh9GaB4TrU8+cTORkLA1+XcgAJgbyjK1r8OSSiSOJZ9pqmNAy
We7Um+Njh4FHMZJk6iXpCKNd+++rHzs4/7ukPGPLDZaoFjj2ccot+IrnVXK3leYYpMLltuj8Kxcf
mcNvwgSv9MRaI6s4ES987M4Sz81TGqify0VtNP/U7KcW+f/UDwFb9m4XR4YVCYTxFYL7w7UE1JRH
KzXXPS+MsPsfnR1dBb4+xzB6CukAd0KWEnVPxswQo06hOvA1cv07FTNbO0kUMVn3PgvqR9ezKzyM
Rog6EaQ/OjlNUpgemjurUqK6BKuWmzCMIMGDX5TRW01ISK2s7CWOwdqwAuepoCyWlEqXr9+9vfGm
olb36bYpYc8B4Yj2rDDxCThVgmgWQi2QqpVVPPCzqQn7KgPTL3ASOH7quIfTaWQnp4tLeI0JVDD/
wasjcPtqNVPrQelek2SD3vuy0fw++yCaqWUcj0UHscuQT7tDrxr4tQoZgkSb8/MzPBByClJymdU9
Gg56HqZnuYtIvD6DLDfs9wDxD5mRSQlIaoax8mQYelHXxQDM3ZUkJ2ea+ZvGX47aL5ljz61o+1oZ
+aRUNASJ6vbCIC2wj9LWQJohteXkm8yClPWfF3t5up445lnf58dnFHPMIJEzUTrohEx/RXeHehg7
6tAS5iLiaB3X8XGs8GR2gvQlAJJTxjfT/xrLOQ2bfvTEvbs22J42BlgnZgps9gGqvoWdKXqn1rvA
Rg6Sm0VTxCNhLY/4n9nkGrg2hKD2jTJWI8/bDqz9Bw95HsU0sgPzOvbluEkAtUXzvvn5dXUbJOyn
GhWatiI3LLeMEdGI5/lFfMtJGMVlqZvfartThIda1mHD6iHSP2mKdpo9c9Pzpcp6s0ZF59giskSz
YvnklQ3QRLRUKrLMfCV3/KSpaOVx5zJaMSPG3zEuE8OsiE1/nE/+hWIxqkOSH+bA1y6laBAcdwNF
csmn0Eh7C/ZFYeRYlIR2dcZoztQnZgd2qvCcPBtbWYXjiB23jw4qBBPMrDaubKflSd5bMSOhm+q2
++FXdU/m99rSKOiXjx+l9IALZfKBB2Ub5VymbxtcaTX19wQ6MCVHtrinM2z5FZJijxhDcqY6vyYT
karfgDMyVjNC2VqVvPTSgXKPbwVa/OmM0xDwlNg6xbUMRcoumAWwjKcZgWIL0teWJGAFtOYTe2lZ
2cNn0y2e1KtCBWiqKGxPpWP6Awg5UihWp7Dhy7L8LOuADxiQ3iEqoYcA04dU0OMUaB/Kj4W2MLs0
ngQiN/IHMxuj3AN8aYMdI6ugnM3V2yBWCH0UbUpBbo0+Al8EyNr3dSF+ITbT7a3YWABPblW3ugNT
nCRKaBcING51cwPT4HpAW2lIVcddOCCpyhqgL5FYiTYCYQE7eKz6j/ILAM07WrhWaspcGBZ5oC8G
VFPXlwdBCS4fPSyzodWaoY2yWjDw9ORw8rgXodvy48qFNgmJMVNIn9cwJ8A7qP4S+2JejGydjC72
fGj9Lx/x58mz77+xjwVPHxoIksq1DKuYxLUd4jRcZbZUSQcwuq4B7IuknzQ9U9ZiJkQJS0ARfAAw
IrBAcmunXWCEo0Zu9Y2cyx4vjSCIL3kAKfEQrZub9CDWca7WtqrN/ukfWNw3h7ql1s9sfiUuAkl/
jL9XQXBZi1p09srQ0xa6y8fwdEdujgAoM4sPX5WQoHyA+BwplIiMu0Yfx6udR0lkYX6P2HW7JgqR
EipkQOm5Hwz1XH6RQA+4Ow7oAtjzXOZf6y4KUb0ipSUWaHseXOruW6h4szCVKrAr71Pd30jbrCuo
OK47LULPq0Iq8QNvsby3MQ9N9HVVdIjCLYnio4lFK/HWG79N3RekM8SDrpINdKH1jxAH8WLbLt0j
CAQt2oK/S9IREzAxSOWFGS9NMSPFAV7FVGfPRbHHlrL4oLxSqeMCb4ZBQY6E6s1dkVZGAolTTn9k
635YsSwaIXx61UxSiorVsfeleajP+2TsnAZ4bym8TVKj92ZblENBBeKK/l2AjrxlbhMh5JOliGVV
d0fsEqAfNNBjUZbyvU07eTvO6XK9R88m4a1mtQ/iPmtO2v/sB8/KgX0aeuZKFqgLF2rmXT5miwB6
DmLzkaIig4yeOdtyYCaWwAtCPCXX0e7UMluFueiNt4+Rdw4JuhMR766Y74Z0NuICHihkKPARFlWl
erumd1eTtkHsgb3XHyjDCYgg34aAEpBOJmAigD6cLCvyBabd+i2UJr/377T7h9qYeJ8IGFKvlO0m
UHIgtyHau+ieJZjQ9ZY+JbImR78PtPGOtjdRPhZquB80IjIBzAAJ2ZxbkHoGIRNVJuyv2LjYXEag
SK1CZ0jhQXiUN7AdzsaDDFbK7gJar6S0yHHBF6YBkb2bQRCdCiFnyJyM5TcOvRgGghO5TPnPrKRq
EZRIjjQfg3/oygjmV6lXEHbVBWcgIMxAop0cmF0//i5qgCZE+Cpku9IQQTAY1KH5/Lh4RiV3V3dX
kZ2kpQ0kQTnG1qqqZmExJy0Z7LY9JihZuTTZc1FxcFnZRsxym2c0Z0AgWb1BDKoupI5YMA8rkSf2
AdM0R0BCFyYCY44C+UfVU5iW9PJOn7aeHR034qW/kT3xKhW2/vEKuMqBupoOABiVq35Ohj+kXnFQ
I0nUNhyYSwHKD43OPYsOzHn/tJFfs39DMRqx7Gsa3cA8w90Z5OY0GnmF0VkzCtLBvrTyuk0ANpWF
0hfnXm8ffqn98PjmUwu2d404tQMWBjxPMFSQwyZEpqWkyPx98Lt8qoop9xd/vuhS1k1COfMIdtQf
8ya/uS7XIIOfSuZynhsp8z/fBgvn+KR+Ygcy+b2OjxqH64OpWAF/95P/2AAMECgws7h427Jd7lWg
8bOiydolDxzQl4L/tRGP9g/M4m9VNpI1EA/ZZf2uZzYRNqxc+D0jJ/DQNCTaIIlqgtzxcTM5d057
Mju0X/kKtec27tPpm3k3DLiM2ngnUl3tYsEm+uFHppgUHO/MwLY4NBdO9YQvo4daGhkb16chTvqe
1t1QanzFCAAlVvpfesiAN0gRrqXIr/CNov3JgbiDav5atY6QTbWlyT4ogCsOepInN4S5Jv0vVdT/
9L2vIU2VZOvGkp2ORzQ1Af00l1460S+TJx1HpJpEzK/D601zRSD4pBV4f8IUHybx5DmPfrHdKpoh
cCTcFnl8GSddeKgc3CPcr+H67/esZG3ZjAWYTBcmH88p+q9OMSrTFP6bZbwC1TeDaVp5td2IOxhR
78Dxpi0SPjqGwwhvg2gic4q8IP27a4E4e5H16mameheZRqJFeZABBFVgRYLh12ApewxRYV3W07SE
Em5Qp3jWp3+MwA9vNMCvpF4PhbhZS/tygRxi6ioIkSsA9TO4OwE8rXmglMSZ/y4vprpUCtaGe66F
MTNHddk4PiNIUdU+2IuaH90Fa4D30Gloa/Pm34mJ1TSyQqo0pBPvRAEIpoKwrPsp6bgnuFBrZVzX
S0/Cznu2ADoTQMjw0l0N2FUoNNyS5Bp0GkLLsMUxYUe1Va5BLCdpOKFIip9c36kGLKhroXVclS2I
NrMd/jzSp6zzmWDKrjDm7CxKrx55V0p0OYJi8uZMxYJq5k98Zsit3S+kQEse257/Wqx7y/GxjVvS
3V4KraET4tJCSd/Ao8YZQdeGm8agX8u5xthiDGPe9qbzyXKSQTd9kB+EMTWvKwPS2+/WHb2PqTGX
wR/ttER5ZfQVNbDU8ATWbDArZBXK0a4wHp5JbNY0UtnaCXv1EhyLdQC1hDIIycNKsbGc1PQ8fRTI
0hJ3j9zxnLeHTvUxPyddvAqO4DLydPeU4iUIWu60tTkPpUpL6RFyLCBFvCcKKbk0nI/2Ocf5Un+t
SAQaip4eRYNW9aXRQ5LuDxmmF2vbdMDFemCSrRVePxRlG3CdIxP8BQvijPCNwv12c/3MJnj2ued2
sFbcY0xR3a+bVqY1/bpVqp72LqZvH3Ldw6Nffl3ALmq//uAEK0P8C/6p5UEtbD1tBMeBLEPOUWYI
qjEJZ7xnvQTKrSH/c8AtZKh1bvhqKLLmhVD0cv1K4GBFVdQIJIQk/L7KieuOi7nzYQ3h0qbOdvpH
D+lTPot8eiC+dpH1SOtul/ul5x+MRAaLQdhKC2EAdjmydCsuIkHbXzswjJCZMxSx6+jH1eyCP0Bj
I/g5ZTLNSjEqQ4A6bNLt+fBYC/RxEsW2AE3oYq/XciExDyPmJSTdFvtw3B5N2p2ts72vc1qtzm8T
PCxsyDYbHbmfEox4TNUkuVTEddxFC4tRCFsPtpvaaz5sV1TCFmbeXyVGy1yW4w7sfBbpz+6kEJHb
ua5UiOKLza9DK382+W7bbmMH0xaoDJ/y198ohm2eTWhPYFTUKyyyvSuvQwFLumEccbGYGCrfIFD0
y430WBo2T6bHahq5dKW7uY4YT9aM8LMvdcrSEv4CbFj0Wwkc3zI5VQWskizJjYETHnlGIMTO9L3g
UhY4DuUwlu8bn0KrUWA5yu9FsU6KNOv23vr8xmmXpW26mbl1Q5VXZPdqZcu8xeY4A5h27Hjm1gZn
H7dj7PWFH+KV4X/Gcuwaw3QuB+BH9Tyu3nLKP2rquZrDCRbVSYe9qGRMn1UVtiTMmXUMuK9Yb+EQ
s1C+foQo2HjbMEwcnbJpR5zyS+WlXSMabWuvmW6fkXBh/WfI+8dTR8AdseualBmpLtOGsnNYJymw
SxRQTFYNNZ01WR1YOX4gFw1R5kh/itvFjGLDEn4p1NrCibS39aaLYw2URrXepLiQ6PIDieMabsXD
dylBcEXyeQ2ZBZicr2nrQhBHgtFfLJE47vdPEa3KeB7tSUCJV8TYD/V3Qvz3GKhUkUsPGhX2qDDA
UiQgdV94PmNDxmNqmX4uShZ3G6L6U/HySeoOMLcNiBNnFDNcYIdHhJnDJ0wLiDkAla0Y/fmj4d9c
E99KUJ0iGDdyflTdysrCcjL+uHo2miT4F7XXiU5ialZc3ydsc0HEXTeZaQXQrZVqEXfSZKbuwWFd
VOit3y42waoW1JOHJ0Xp3S3FoPsL4HOAkHmhsEFemplw32HOhFrGpvEDdmef85R6ojn3enWPcq/B
s+2T+mZC6DsYN8t5wXP84DFV9TzqJ/zimh/h+D+7zx8Cz6UwFgOIpNNIFIw9Sqo39FXd8oBkQwmF
nwnY+I2DvyrWZpPnSJPD5YwSHnK3mzV6pS4oVzvqODaOvbIogmAk3LKxaStZU45En7Uo50s6/8fL
txWtW1V76puOx4poCMsztXZoN9YoplK1v9NEyE6VToHvgAVgi3dVaueKREISHwwgaPVtFy0IJs0A
H0Ofluw0ER5sZYr4ffPds5TWVKRMzLz7y1R2F8/8n6FmpAAwKubSjSW2BZQXnFWF2kCplBcmqExc
1hHO931c3WatfAV9N2QBJbO/Q6qmi6eokiUYhFT5fnHqJQSKYjdn5QeL7TCbqZpVrzPSsyY2a3PR
309Gh4OMktL1JKxUGNL25qUIlLydg0hxS87xm1QyePer90TggirFaqE4fS9NJ2qVet2s7y1XRIGQ
1Lj27oSa5H9h5KEAmw+YElcqaymRL6bm2+flhrGYrKa8eYtbONc7ashzCPnM3Id4oHrQkUOub0D1
2IGK1WHgz8nPy/3bBiUbWNijnhOiqy1tF15DnZ6zDTGnhbzHLIQ0NPgH8woYVCR0sIJe02WagGwW
VEzFwH0FIV1AHu/F9O+5wRh6tgBRQouHPO5ZXON1S4p4tuBxSjB3tI/61e4takdX1K1c/SZ8Aysf
fGtFgGTXGWs6l61s43p0DSwfbWQmA+sJzZGB9RssXW76NlkxwWF1sR8M7Qbiso3u1qr/BIsr+6F2
jxNgF9RQYKTJMm1AhemBWn/Sh8XGjNQUQK9j36kfad5o3cQ5DaEuMcjos5Jp/73xzduuavzq6u+x
Lhsx+KfStttBh7AbJwJrALnNmdqg88PsB4m/DF/9BHJTMG4+ysqplYjMkh54Og6oZCc2/Nnq/txz
0PfXAWlT8g0vvImLlEdwL2dHVNj9jO9AIi80ghpom72BLBK6K9x4a19uv4mq2jDOPYjy4rPLsadB
Q7lL3SbX5TPMYwX7h59M20ccTGcfC+C/EMfym8XeZ0a8AOdHL3G+XvdxPTlN1S0amgCTLfT2lp6J
fOKXnAbJLCRjmw3F8J4ZHl8dgfJCzjuVt1yitfbs/Vbjg0GBkNUHnK08efble7uR8s/brxGbrjKC
FNvV2/QTw/4uz8AbNBmy6mfjvKrR4GMQgXkmT/gJWJGJjiOWfCdeE+fEhhS1EIsI4z06W5IfPJ1i
YIccx1e+H+YZ4kTAq9Sdp5PVwg9/bUdNJBI42jqHlOZzZFcMYuQbYhMrdvv4NKm+PpeBEJvCcxTr
H938/xuh7CPbq9iUP5UZfYpCD+tz2QNCIb0EOLjZ5RLaLKXRjVJpxa8doMgJe55xiQLTahwXQZvn
AXsj68Fv9RGGQsQiXqikHJFOt4EDKLJL4p96I7JrFzN0H2vkINNwIkca3SCYl7rPj8PCliW78OLT
XCpZBeSJqDP2BPJqwOgoX+F7t8O8OdgMsonCEKlglXxO3OuedLYVEOPTUPWHkUqRM4frUk6f+nZG
tqYP4jC0Vt2prxfyeBHWxly/u3daLmds/Ilm9EBo2HPDOmcx7hz++PkSoTQsVXkspDD+uY6fsRTc
JPyhKUVmC2PvTB/REbjA+HbPhFuk1ibBUl/P3mhrUG/m71Zb6+EODSMHUvzmItcP6ZmxhnWljKdm
vFJBQHNH5hXblCYut60Vt2mQjDe8pN/h8BGqbZPRWcTXWHZkP00sb1CbqvP70qOOpwysAg8sFQY/
SIfgp1DpwUuHxqsC48ZJms0ak+S6SFrDpE+2dVQhs7Qo0T3JmoOVkyp4CwCoEp8tQoC/72W+a9t6
M2IXmkOj2fQl4mOq1Ftqh3AvdLkQXYHHAG8rOnjpZBiYZhw5j1eq+oG9nn1/4cKjoDVbz5H3tt0E
J9zlwhnV74XpgsZ03Y6A35qhuBM+o4VPNMGtZt9LMiQULmwM8mPxXwLo8Fqq/CpUP7ejb7L5FC+8
9r8K+b8fsCU6U45cAsBdOFOO9GHhCFXM79SXaRTMxoPVPJZGEPLP/4tQ6uY8bRmUj1zjJB+pqut1
89Ns681PBgkkpjDzxjDiVfD4cePTMhCJ8v2r4/8hqJWt5RAZzYsXpOLufBFzQz33pjvTZYahxNb7
6LEbNhKdE0hMM17o6UCdrHBrkQJpTZs1rdriyspoSiLRPuxTEDJ/mwGzMZCvEoeveJMV7zcXhtPN
2hha3cKEHVqBgjdAhKlq3OHi3+iwsfaPSBpOfeh8+Y7dXfe56HIbABaXeQ6optX5ZhqObSyBNx/O
kYn6Ja6d4WH82j2HZoMHOjpE2m9Lmpmzi0STqVY6nmdLJooN1ohz7ZrTCLCWO1VclEUn0hf9sGNH
/v+iJpLlSdekQd3eLjAtfgHhmXcvrZ/ArMzOit9x5Bh/X9CdJwA7e4mFoGtKGtvJO2et+cBVeuQg
HxJ3GOWE+KO+iT6/FsVscNYN80cekq+Mfe3IXBXQ037ZU9eQiXoPhvKhlHMtZ9cesJ628DioukrV
AImD07SAn5SssZgPZ3sGlj/rZ7VKQnElK1AfPzfxM+Y8mV9tnm4mJjzHs4OPDmv+HhPX/oybomXU
t4Wbe9vHZoQrBHOWXKT0G1tCfk95yMpjCNaKYooKklpeWMeQPbfj7Dbu+opZVg2l17mmUkcs6Ata
aysrM5DuE/XpCmeugpM9LGzyY/rQBaLsV1H9FgYB8a0osQRFwFhqvyz/7s/Xf2GngQsObVgtt1HS
1Q1dX5Z1K2XouIE/TfFbMyHlvBMdx1kJfU1QeaTOqzABc3jnPEA507rJ2OUTyAKNDpCmkS/mU5Kw
flj19YFnH4b6baH61uRTxor4o+mfL75KGdvHxc30/EfVKuj+guRRYBxKWAcGWdzCZrja/6lTTvj8
lGck8W1umlQdCxQ03ECrrhmxwD1b/lML+mQEMryU5+tF1bQkkATKuCy7jN0XxS57z291j0pHUy1y
iSY11qYB9SuEXvlVcUt5aokzQ7Isplupj0AFI0CvoHMYA8oRSEJbmGK1wXljYYXqieiHBiBTAVq4
cDqWdu5RoCRE6HJcDtM21cvsvVED+EEo7OvDKpP4v4ysgJsh6In3RQZEYeESsYvbn7ZsybpUqjVt
UW9J4Rs9aL9t06hcPBaLUtTvAmJMACbX4LvpjN4tsOHsqsHjjrLmJ55KApRYP0Mv0Gcjn0+Uo6dy
ymI9lYQ072svjiMK1ElxmtRnZbmXouIDVl1pR5pUCEIYSqgxPq0iuUGfoHLqSmxe6KgA4sZCzGGg
HHkIc9Sm05Xyhq1IUMCa9fwzw6CnIVNK5WBOqzJ9zpgE1eMT8k3HeGS+ZDLIMI9jOTbR0EgPo0+W
plOTLE3qc330M7bjgmJFl/g4kfFbqG3Y6JakkY9Mz2DEP7Ta80lkyU6IaI1bQMtMT78XtTFBave3
mBzDFYV011zWywEIXuVXWhLzUNVlv5Zn7aXYrimr6lWWLCeN4wdfqRnnx0XwhDnWcSXBX7FFrlt9
9ZAn+wm2OADn0PJJdOfWT5wNscE/GHnbd1y0AKDce3fQdqEhk1lod0uxgifhyyeAFwq+JyqAtlpb
XFLFcpRlbEwFslQVloKTyD93sHkr4a3SYy8PC73LyL+92ssOtAgMHk6wB5fj2xohNcbjwiTPHhzk
Q5WO5lEH5UMuAZhN2ihvoGqUCfc6FFCDBr2YKJd35mOj8L6EULaNpMla0ExOSNESrgBJoD+62hT8
h3A4mV9rB7zTKBg//+UTzUwEokWXw2vbe3qablak6z75BQojfDE2j5JBAEOUPM7YGqvz2++HknVl
GarqqkVwJ+J6hQX2Qz//bMubMwZsX7LP049+Dx36qewK9UkfOb1c5nSINkc+FYHa+V81aWO1ryPC
uAxtBh6esNYZK3x7sEG3V/sk1LDVD/vDUFLBMu1pUlEuKFJqbgiTew1ZWL0RlowJwbjJm8xZf+NG
QTRQN8KwIKVe6vP8q3tx243aumk54ec/wQBpaiklI+cYSfWZbey+U27/UR5NebLjbRKk09iRxRUm
Xk1do4xzHvg9ld0hArI4eLZ/H/ks2M+Suh55yp5Tq2PY86iUul6rrzC2acfTgXpNNbYEDlGn6GpQ
P5GhDv026dDmspbrVP0w6y3i9toHv5WoMhMOBwjiUBY/cIK8fFmt062SGl0AZwhAz594TT8kFZ1y
moMvqtK8kthjfkAv2m3yAd9r2qvXBc6APTKnsZQQBzcu6iJ8x7Y0M8w4CmlK0AriZ22yn3zWt6hy
HH7Pj6qOuSzb3gecSq6sgb7B2Btsd7anxajw++xuSk3DcqN9+5w1Qwpp01S0xB3W+bs+ZH19LqF7
oNs0n33amYZVqcb0J4//Vo0bEu2vqBUROmXtMzBMDIiEU8tQ+DT6P54RhG36+62GtQZ87N2t4/VJ
DKtnjglEdqxY8nSdZ7qhkKCdsLkydP85GOa6ue9Xa4aoLIGYX8EeoOBsCAzVEkY9Go1jsji2WDZr
iYdkh5SEiTuJth0ZYiup1/FlxjFlTgKpo4Ir9VMqVXFutCwoWZuNnD2eZgXO/2t/foOsDSQWKJSN
bAms3U6W+JAGFzFA9K5aGAV9zbzxrp7PmDl/dwCumJTXvGLj0uVyFjBqiJwRGisxCnskky4gu+pU
GQZZb0827LzWKU+Ae2xcVtsCXkzz1zaPaLx+62XMCdcXNuc9U+la1KwX10CUasOAu5Wbz8M4MlXY
NvhHNyd42+8pTqpglPRIMRvbHirssT8Zt6qlssad3k3Y2zkVk+9b1sLeenRHrBd+UTOImuHfuMdz
BStpLEaglvvw9QCWAHEZhAQbQV3FWVRxqP4QYDbH+Zxw75D3+nOXCUVV4C90jNkC9dOnWZxyEVfb
vHrn7PQU4KeHI1JqVpuE4OJDqulRxT3UZi8YB2MW74fgfk9uGapobTWyBOBDBR5mIAUVSts8VSLO
xbNMMLoO2Phs4TsKaoeNTLAM7uKhyRV2ChZ2CORBfsO1tZ+ta12PSM3AV1QJpIgpP1YqtIxNG8SC
Q34uY2p/8uLfc4m0x1GOZEXg+I7RwN2b5mKxW8dFoaKKjkNIvKcwr5KrvEVRVhQcTG9MM8KtDGXq
2MDk8XgulZgsCdBC3RoH0/TMzAbnUfZKUfjuIESKWOgd+r4T4JlUVD2So4xMD6KtI2zniqMvGSyN
4GJeNEgJ0clRlv+tqSKN9PWdo85SGmF6aWu7QsL2uEPO/Yhz3Ue0mtNxoL1fqyFCbohYCGnp2IG/
I+Rqzt6ZaKZC0G6xi2mvw4LTTIBjCOgYhi5WmYnwIPAIIMo5rQVptInFj9rcHaeXDnHSP7vC82vF
WNjVkXqMUxF/PcYeHmA+ywe77rYMM2eArFx8MZI6zbPnf7YmLBhApWdh+VcziX0FQf77jbfod8/J
TqEDGcmjehI1fwUoLXMCeSURkAM9ajvsX4MSDc0VpcmJMiw7m5I0VOUFEU+J35k/7hNQvhdRTYbj
aXcV5UzZdxc6cbWk/fobr70VpkiBvTEDOgOzssJ4btf6mabbiYYjRjByJgnz/vnirGvT0klagT15
0sHXtfEW+nARIH9JWLHsBQAFwB0e/jXzrG55ccGmGQVPhQQsiMxuttnKFJr+pC7AnlFiarfnVfBa
3ROIwcr8JVfhkwtpiv0Xq2PtRB1icXsQZ/5lcChF6HPLoys2pKgQhYX830+wBCRBRwHXGNHaGL9e
W0mWp8ogqHV/nJifn63GG4/l3gQ/PQHAL+xg7m+X0HpkzDKDEYJgdjkMJXUmfpn72cHnSHEs1VC+
JoHsifcUrks+bAgSU8rkOfB4DSXPC7Qdg2jCt7AtaXRLRgL6GTEPF7YdUhvJhFgbfIIPuGiLsi6v
4ohagUbFQo+G0TBz6qG7BVZuNL4OiTHIcFrsE88p0szSBRoc9afHwda25b3Y5ETBDlXBRIlIFa6/
ez26hxb48Wm75lw7/o/ctv94+7H3aKYqyp8FCXxzWM4E1M/VGXp4zSm1EThYOv6icGO+PGXIG5ar
9Y9jDrx1wWApKBrC0wcA4GCHcxMwsr0Ta8d5TUFeLRMo3x4HNRoEI5btgsUoq2rXc9D/+7Drjdpz
FRVsncmGj+xeOMxb+AmZPgIqPara4ArytsqdSiu9dwJarbS6eEaNvgFpoPNNoshUsMBiYpiBz3iA
JDAOzs91wNLGELSgNIfFVMBtX6iqMqroeKNJpst7b5Saeu0zoS8nWcJN+Qayx0frh7VM4cV3gG41
mT8hoKSz5mrP3s3sJSlGsX7E0ZWL/3nCvedZmvzTkzCqcLHDww/EzWYIqIPNQqjY4YiL0NESgj93
GeJafNrGGSZzYfoaAeplvHX0t+SI2P466Mq3yJEZOCwmC4SuiAHQYr35K+MgJRU+olcx3YIsLVpk
QM4g5Yc3kPHP7blMxtBPbsn85lf0JLCXDc41+h9SY4a2jhsk/7ENKg/wC1Btn4582oP5XTIlP1du
5qQoEDk2moN1Nx/VENdRwx+TcQCLKjc3wygT3uNmT6g1RsEWckfAgYlqTm2p/umParLRkfOpUPB2
vGe0iwk4pkvbFwKrHAwd9mFdbNxmJzDF2t0aT7lmLMfWtORPsqNjGLKeUcDzPiCF62xxoVPWQ6bg
59v8dQwJOP0eLSlSYUouYOfBwIkV/aUo7icZ1y7RHTfes3V+aKj083weudFM3CTYynJ03SXGuHt9
EQdCFkh7xoaFm8yIv2S8K+HEM/JiBzlyH8KiqzcXk9BgjuFfUiPyYoZhBk65PgM3/aGKZZgDFHCT
1v25e6Zh27WxxXK9NBIT/3cpUZS5lUPdImd2xxUHKvlnxsrMKStIdmvOkZrmGIQSQaz1Sl90nUxo
NmY9mOKNrVWKXMEBzNGeG4HhrQ6wygGjQms7yCi8P6Jref+CgkkQfDsvSNSDuySUq5e29edjx+Kg
OHjAbhHg/aFX1WTeslFpQvp61/Hdvlm1VIWUkACGPSyv7DxkAWORzBg+0L6itrh79d+aR5rzEs6d
BLRy+vjMegOMcnNOE9xiL68j+UwsJYdS/TI3WjMK5F1lA2vKpagx0lV7ji5CzYPX/sBZ5atpCXyf
RVNtAwDsBJwJj4OAXp1ydysno+2dJ0VHItt3nmfLWHW9khE4npUDX00hS0wkBFb7BSZD51Tqlga+
8P9/NAHVdY640NcxBE7A9M5N7uIA+MkS5P7qgj4K46E6JzePDeFPitWWw+sidGLfxwkjm7Q+Fb/a
j61jw3RdeTiV+1RIpPGUAOyWxzqIf3DX6NgDryGuh0Lkse1ZVikth4cFR6a+fTQqH8/CIjLS83f1
oPSchjzhDChhMOI0WWhsyqpNz7o3952XowzaFLJI8rEuaKPGXQxyKJ6lA8TAsVEwHzNmLba+gI5i
agSQ2PFh8/Boz6TBiADf8cpvOSAn4SlfjCA08RZybWSi6nvxKtwMUl5hEzzqhgkB8mg3xF1z5g0b
xkssaOIJ5Jv5KkFu71gAKWCNowe9e2/KreioUf234jr6uCKuSQYPBhr7/8+OxT6WBBUNNVr1pjF3
ymPSWYNtF+BBik3z1NqerDQGmSRLJmmQlqxT8fhG/a59sMfOTC/zUxS9mXTYUtr4b9k4idbxe+hK
VMH7gEmc3j95+IMYMOTjsJ0mw2HWYySk+QL4RMOLxtNWUSXD8+thpJXKy6diiCSc2qsJesgBIKVL
+8CxamKJLu9wOyA/o+Cl2Ct4aOzdMwtX2yn0cqB7qhxbjeD+HlprLGt63K4Hb9/t3nkOrEjZv6NZ
zYU8OaiVVOt6ddsFijs/S1/yv/lWODbXEXUL2i88b22SaR1K6RjJCLPG8uXmobEZ1mdPFPLkyLLw
agYaaCJcbZIRwLJO8WIAqALXumDkz8iSiP4zOVGQNHE5vBJgMXH9q1k6Mx8K2ZJVA0fjm2eFM6il
hn9VtMaWjy6uu1RmgLWUKhEJpFFfg0E++MTrSrcUm45QuyBsQgwg0ai0xj98Z0nF9Hud595VyVp1
QGrK229tX6Nw1su8cAhcxv717smxlZ8IxEunVfOPRsns4JDW/QOrLaJr5Bud4F3TFaSs1dsuYdy6
F9RoMyNIUtFR/Vvrj1HbVMncF5ZLYOUTrGTwafmJeS8YFa4HB1fwGHUU3K8TFvYQZ1mamVBP5ODm
f2DYrwjSGIO19wefmWM0IsDZWUOi+5c7Hj0K4sp6kQt0JWVxYMu/nvbOqs2MY793gy6/jfZPFatZ
r/EtLsvLOfyU6ODZSOTl2XCuFYBjHmSpMp74VOcdinU94ZlN/xBhCPhX2/0oPqDnpyAouwasyhYp
KpcnnXUvbJHum5RU3qmjomO0mkjkh/vc9heNoZTUnX+0LqcQ+mFGtXm9dDoBeUFpGl47CcYa6kEw
NAnfhCU9MBMJv7p3ah3vDWlNg4uMRLF3fxqUiI5wkzgyRREBRYLXn8KsTX5ZclM74JrpqvETHIKX
Vv1bdBXnDgAKt8LCtatJoQJkTUOTkcq78U7PwIPk/TjHwpnAhRcpYoHwWtIAfbEOmYbs9vrzk6VT
MZzF68OrC8KRJqiysNfbjkjI1GLEFREXoKUVC8stqT2aFwVvFqEz4ZhoBOl9dnBECLWjFl+ayiLa
KztUumLwq/ChxOEne2aQ9qbMrt4C3KXwe2p7ruEJ0xuIV3YgOXQ/uKVgXS5ZavbqUiLmCKijRRbn
AGTU4E6GVsjMVognNPOy7DgpHS3gok0q/v77b7oA8+W+Dcp84OD+FWkv1ljaSnoVJIWleBQEUCwq
WcEzne2daOtTk67drwZyhIlDi/uCThwUVoe2HMBdAiaZBJdAqkn5e4aH371/0PBBUWP60eARoXnz
6M7S1eguNyiUvvw8ZYVvWmCEFyVl9NMIM5B0xBqSZG944w48q0oZICmOgUz4mKQ+xvSYARzILOrl
PSxCj3oDV+DH1rzTN8fmAM/ZlLE5VaqLqNB1uNLZYm+qTJXmKEOWaxSoN7SUw6eNd6p+ZJdwoam6
x3f8oLgxtMsn9wGSEvP0MXmTNSNPTh+cKLnHrX5xOKe9cKWg2ANX90vTqqxTE6osYXazZT+tB0+r
1GmKrLLGDjn2/pAWie6Ge6iBM4svFxs6sqo9tIkvU7mBhRGGrAoujrE4Hy/tAMhCRVuVU1iCrZm5
WhP5M8iBzrsRG6/vNC17BUcWTQ6cjZvI8NobRlRwIghPXQ08SAbgBwIxUHXehTFmcteev92f9IGu
Z9i9s/YrxCAO4/aw5+319LNiTS0qCf68T8Xhq9X4jQC30b1OISQ+jjMcEL6tHKz1gA3cqPclIwXp
f0HFp1FCX17OuS2Q7yTeFktq6K+8i8peI0NqAxtLN+F+4RstlK1z4Ha+nkpQorVQ2PJ4SW4N22gK
m/OTWwR7q8Yse4Cyd5+l5RyLL9SxVropE49cKyPW8BoR5UTjvuceJYQ1NE1DernO28fDwT5OETjL
TdqQuuOYtMLmteSw70r2s1sdviOgmrlqvzQ4GG1AQ+dhnBgIEtiYTMvoA23vCotAzPXCeMyLrXaE
T/AQEN3dm6Sq/PIbNy6x18Y8qF+lPp8+YWcn3ky3Ix6NCGOgkH8YCCGlwiJGunY4dZxoLKlIKC1k
UvwMlLi7PHdK5zmXxz2jZcaKWXOK2h32UaThW8H59BB1Ju3YRcmtwfUHk7fRDnB7+FFYm+hwcYyF
46h0tod1L60bLi+jt23tbzBR61BXrDQbHev5fZU9FDopyW9zZwr48VA9XCs5iaB9yNHOfxDR1e4y
axev79c3Ktz7qtgAOmL8DWpYWiElRCMzXtPRXlUMlHPFBj3/TsvkNt/B1BaShI9251jHG1hI9Blu
dLL3rkH5Sx1Ci/DQMQehpE7Kys4GOCsY/hWnnCADxO7dff9CV/wTSsMyvZ6xdZeGYeHhsPll5E/h
926asPuSGNE2CLLmG2UorkyXgDf66iNYgIUK68Fht+FLupBDhSlggU3lPXu4W5IpyyuKLQxalqBH
jVy2StHdDu3M0gD1vUwn68TqemI8pCAU18nQRGm1LemBnyWtphj8n7oFnHTjpcwjLwzZyw39ZkAN
bHO5psHs5ZO+ZgNWtGzeJNX5v0SRtIdBgaDYVRdx6fBXmWZ44KusTDBUYg9tkvD0pZxg0k6XkCY0
hnJDQkRpUwTjGfkmMdxRy0Z5Zx2c8tyVXeF86JNdZY0iw/9CVM0Mj9CjvAawmqc8+/qcT+aCd6IG
/hvf2SkHU/uztVusH04xSHf7YLmvodij1ABtO894mZmeM03p5GY9cvOy1SgRJ2voUzdREvM2i6XO
xdoYQIkrEW2cj0GKAyyaokZ/0G2SshnH9Dm8euoDrbFgLLrP7I4ytUj1NKoCaSSTV4WfmqgbW7JO
D4Chs0Nh8IMu3tI1x9GdsuqjAYuqUNt5yKLWhKn3rlvkUZawb13pR2HeHMhc2uZyy9nqZEOWmla3
zjRDJ9tRD2wqgw7M8M9jxshvM8AbuOISDyvqU3P3DFGuHkhY6e8DX4RsAvtvr6SC7DDx7QYu3CRY
cxxmdPh/vUAUkMz/YF1MDWiwe2NCiNwqXjZ2i4tlOADNsrOX3bBrKVKWTF9o4N+jv+/KP/X8WA1e
Dm2OE1iihK7Qk/8/436R0fW6B2s98+v4ZN3gam6t7GfEcxXc1Nz+7IEKhKOOJoOmLDu6IUiE+iiq
Fm7F/yT8Q4ueqgPbYnW5yfNowHXIZm7QiG63PQX5/kPQh/5CpA3XxEbXpZPMh+bY7y8TJSIeUdUn
+Alh2/ABjCKyvTPVCQWmIAeyKO6/iOwIwyQ+3655N1Zooic/2oZaF73dKobEc5F00o0YmtXv+P8/
JN7kTDyKgh0/HjYnlj3JiCoZk3nEC0vxq0csAU7hGOjnMnsP70xPeBtVpWUf7JOfmOCwDBSqlLZQ
+7fr7KyoBVn8u1OnsR0BeSoHeapXQjVNtEXLVKOmrzu/lndwsTncw0aIPnPJhgmSpaTBeKzEO+b0
B2UaF92IXwNLLrOpDyuAwz9w2gEQOPqC+w0INu9S/LMU48OcUsybNWc7OHT7mSpA5vLXbwpPdAQX
ySppo0hHG2U0H+pT0ri1hzcyC3xf+94Yi4Pfz9S5AxHqtM7YFD7HnAPvV/lfYJIF2hnPpMqOniNF
y2SlY/l3wWqayY5eKJr1E/3/pYf/PQ3RoKbxSQZTy8IE32ZXkUKpirwFd8U4PVoydbrDooACrj87
8q7ZC4yqlDIRUcgL76mePX4ZpS+DVqdcZrNEzPj5iE+JiiVo+Ui5jsdj04B1rN18FX1lUEF9n8Eh
WdKnnL8D8w+uGWAp+ehYEDNiB7licKw4ZXqriE/FS6NEj15fpCj0q5WKG+2pBzQwvx1taZt7F15E
peg+ZGGU+OIGL4eejlfzodyDiv0k//GfKclGtGucbSRYaIeVOrtOxbCLkOhb+VPZj/nqQVCNJl0S
ewXTKcBs8Mm7zUPImgF7iwVXDeVnL47AxDQB38dKqWN1qVojs41Eq/42Vt/qBixgDNP4XMubcPKs
6hUijMOdnguzK5jt7X9dH6e+1PWGuJD+rj40JVzqPaPN5FljZK432F7m4Ta6sxLjm/u9T9791wdX
PF9PiQKkvYn8USyB8P2POO0NTn1BFo6vU4h27WCOCuvxlz/bcDPwMTqnkaJJwCQC1PZIUukQa5oK
hhulDA91fGcHk9L19imtvyFfgUtd1l+VZRUlw8L+mFrXIvzVoXzr88lM+htJPtXISwTDFHL/5AGn
bCm//VAz9eNs074KCW9h4jMu4CFxSqgcnMVauUckt6hp7m1Nw94QqfkMzTVRIAPC5fHikH2bSSJO
/NDeMHv0Su/263s1DbcKTpbkPDkPzdxo8KaNivaF1LJGfJU1emXGoSs56LH8ON3p/x2f/o0xHII4
NTbK/uWwU1J5to2ctT/3vNUxS3SxUTxgiNBbqjJt4z0rEvdbJb1VJ5GsmwtRUVGr5EzJjx6UDZxk
wt0BkNT2xDuewv8iHao08ZaAtWaAc33zPlnVSCW65DISdeW0kVMtpC4NB84cEBHwUWSee/omSYVc
11DzIvADQDsvJIW3GjRCPW1hSPiLbHsAuJ13bNTlYWRA7nU0hCmOvFlD4nM9hwmFIllaIcOYscdq
ZajjPEl0qVB7L9GxX0/eq9k3PNhPmFhzkZKQDCbYsk84hA2wqMkU/hK+dZyNohrZdJMtAk6DFhW9
gyxgpYiLeGNr0Bv0FrKwdEKcy2ViMWZxPVYeFsEtbsGMSJSJISbrSZlrgzFBEGl8f+mRXLrdDLis
Ps+unD6JU2K1vpS6RsLiE2RA7xLj3p090wPs82ApTKLr4/+iS2fX7bLenAGlrcHIu4cITODK8EOT
zsrHsiary4XwMKJhO2xn+MzGv/5L+TmF/ef7xgKgjS2KcbNMBCn5gPxT3PWfrx7t/2HW4d6ZDp5P
mh3pJm4KzxKOv4k6/NEDbCp3JD+/DpxFzn2jsgvJEcASMu8Wn1M27XAuLfNya3pMKsmyu1sDyICD
FC0C9LAQ9jrCL2M0xEo/D1r5gfD06Q0/4CJKeIzvt9OH6kMQQTda6XJMB5gy2TxsSwnQM2zP840e
nIYrue4CRFKuASZMPZSmHupudXjgj0aDfiM5T8bdc8NRvWNvHYwUxvBCm+cpdPNuKz4Oh/uqiAEL
iTiTWydn+DG3p7xAkHcm64qg/Ic/GigF1LENS9M6SttROd9oQNJCop2qJDNcjUK9MS1SedzbV/YH
m30qtykk3sf2gur1AaQP8i2cFuV8a4lubNNNhryPBzv9BYa9/7aWBlxtv8WapBZsGeEEbERi43oG
qrnpEHGH9CR++195ROHNuVVLr5uADS2gLe1XheO1ahSIufcIOeMrC/GbhrGJ07FCIwtDnQH6mBHW
1UrvYfNoY4UQj+afpC8HE2diXSloK20MqpK3B7mzf+xveVI/WuXsks0DUrypD2/hPaEGGHEJQwaK
EiBozflqWtKA3VOxNsVSEoWSCtTnTFj5naDEs5okyHyR23nMzVYD37ItDPPpO5tU3y70OabOfxhC
V5SCtfj8E0GG9kNR+Ov5Arw/+KOydC4VIp4NQ/MwR7+SuNvmODEjPyKPIExkZ+G/PoK1Ew3i3/rL
bowZeyCzqzd/PfXGKWoWAaz5w5P2I8PO9ByLCvG0KK/Y4wFsdTcgCT2/KrcfxhxI7sFDQVzR1Fx5
ovJd5WtnWw+VMkuPyh9Wq5LwUtpffWT3mawskV25yQ2YNRQq/5H1mrVV7r2miT4lYkcWLNToYKvr
GHsvzzTSPmYer3M6KJDkltiZTNTBIhR/Dt5Z+mRcxd3j+/Udof8Ek/cAnzfA/zC6R4Bf9qF+7k5p
VfN1yfIqUenD8rHG0CJcl+UXNoddpniw+258JFClTjJ4xMv2h81YjhxpHUEvTb81vsnWFgdKNxLa
4HWQkl+0qpbEpGshtf0X2C9JV72IZ1XFkGUqDYbFtOh4itEKpU7sSMcunSg+QJIVvf/WUuZOV+wY
bxrxN/Vq52Np/+2QKAtOllXTbnQ08hwnPlCoz2aX5hDMKaHRp2ZZkfKroJ9N5XvkYElE8MzyO+NP
8EmI1eGzuyxgdJUKuic8oKct8Z+iIEZsO3lzd+7fZt9E3M1/wX+xr7WfWxnG4QSaMr0Lts71zl6U
8rlDVkRM2FgnVYr73bBXnGyiCYCmgZM94lZoodTyJQWhWiJVXoawvNZmdjJCjH0iqX1uynac47se
jyl0mc/EfO3/+yXPl4RAcPuuR235RYm4P0ugJ7NygCBGQfpgTBbpXW8wTZ2J9sM6nUxB5UHbkWYP
v6q6CvnmN3YA7Rw+3Objg/RLZlZAXRNhN2j2CO1snilOaQJZq02k72kS3IcIw9EgelwP8HBvvY0E
Fp5JHpG3WMRckCVu1sc7BK18ZYgHIulvWlXL3JpO7H9DZXBuhPOZRmJdwJHS+4IH+u6TdVvvHyb6
4e1gJZ2xa63BwDOSkvv9nRcaq4ihufGvsIaTRT8aB3nXE7w5w/mFBu6k+F5t7ysyurSwtWxmIDHl
7hgbILp7PB/6+y7NQc6pDL8y77qpuQE2w5KWHzLbkJt6NIG1iWJDVnTXHt94QVadd+xIuXQRKZ3n
Tr0bn6wjuJI6d/YgsHm9geoayb59m536+a/bNLDDXUKLoNTD2H6u+R0su1yo/frh4eyEA+bxRXax
IfAabZ+ZQ38I+XVr8vhNCg/Rwzphnb/L2X7M7XlACxDNK6d6Oon/FFwwgTWhgIlXPT+n/neJOO3b
KsKxxQ2ykZGPJK6HZcUQ/axtWviJtgf9OZS0H4lxY70ynGp1Llg21GYfOIK2Zbh8LxSgOa/2VcvE
2+B3Kg3Ksgb8FGVNKLFH+llpz9gspFL2PJERlTNerf2bVD9ivwbL0ZCRox9OtZI+Rhx/bZO1ElTi
0FgThym+fjfsTvteROtP19CAdWNn4msQ63iDo9pWcxsiu0E7C1Ykdpk5UTQj2fOkYT4qrBbVWxwG
zNlLqpQ6Rth6h9aUFHQYofulY1I7q5k5oxNlZ3XOiy3MOQKT46Ff89/1lRxEWP3QmuiaCImLABj0
QXhFRtz42JS28D+muR9EuK5wTJvgL7z3JGt19Vzb2uaUPRv7YALNeM8i5sLTLB7MBw8oLDWvymlr
8TwYD83Xoz+LVQEDStC1gqx8rbm7rMVYduUoMGm/sYycl910WpZJQ2tS4KX6TM8Cd3VonOB05kbE
9fx7h0ghiRr+ggnsbefiqnkKU/RRUcooa3Ms0azLYBRClocOnRlQJvjLut7YD5aavVEMtHqeNFPD
/lGLMqJu4x01IPRpSa6EKxLHB2eEiK8na0I7LYg+FCzXS1/xabwUCYIDpFqaOweGfk8XMSoCnF9E
In20uTakPuvdC5uqN3+FLsGyXotPYGkJXeyJDahImHa17mvK7rJH1UNTnihjp0HEmyEAAuhC2A0S
NSgDPPigvJDH5L7aBMJFGsUd178YbsqiDodSv/jkQuo1McztlRFsyIayM7mVdiUFOsV5EOCDpKSe
HFbX7llOojK1gLJ9eOwpGqHUOnHMa88J3oLTytjroH5zji866GbjlSmdcjigmF+g8E8P0je11n+W
abS+cF+KL0ct4ouT6nf6E3nU/MaYEcbCFh7AMDa/quVVKGhWx7VrFXbwLZCn2NnK3szKb8d+SNIT
RUETSe0Q+kQagdhN8Mue9e9DWTL0aLhHmSfrlmmqzwoQ11N5tOD2zOR0L6Cvqo+QvBrrw197UQzP
C0uv1SuWtZxRalJut7/Sew5h/YBt0Dn55cNXrfJJLkPa9HPcmGVVpfXdx4NlfJpc67D26qWrw8sL
wuRZ0HfI4V+qWt5M9Sc66pH9Lsg8iQBYCFmA57X1H36KLO7w9dtCjF4E4rWG/fSLaKftQCZq3eEn
346oFhvFeXCcom2ehpmXHKtj9Fc3ef2uvO0rI+BLS7XnAh0zLjHDrH01wMgCfBRaLlQlaRTkV0lC
VJfo50NPRpTH+LxtO1kHw5e5se9Q/dumQAnEbFJPhAgOmSeom0zlNmxGMYV0ObG5ZeuO4/8E46oj
iCMlIDblOEvxrRYNPUD86klnscyaiJ0nVz5f1gio27pFPDVfkhPIvmoZO6bkM9iy2xGTQWygIIg1
4QrE3qmqJ19a05mqVJvt6YQYZZiszbq0gs4TwQTOqUesGJ/u6f3uYXCMGVGTw9yNGS18vv+Y/jlS
38klggdJPfkzYzNo9WvtgXJCOlVqCIvcu3PBKpca6w3PVjh96Z/iQxtxawRUtVoGwe1mYWHf8ExW
Px92Gly+BJoaHLua9H267dn7XRlhLW0Zx8CRMXL2UqYerbG5kPGtglsINGzNE3pDWlBkqkHqE+ZL
hsAJGjxl1rKbXM0Ym99BNp6lQEeSAzZvHyD6jAa+6vKqQccwCKn96eEE5NBQNrbG/8NG5D5fGqmL
1VjtJYbpDThwXYW5PGFgT4NuEbpsUq0Romn8qZ5RIGKyyMidjmIODRFVUF1gMv16ktA6W9NvLiVq
iNgjlV565TN5V5vUhYcCFH/24n0GjN7arOvKalRULQDgK2NELnI9JOyOSytNNSbzj3XFthn99hn8
KtZq3g3FwYd44kXb+B4mWpgPakFwSO/Xl8qkM+jEVqTRZDhhcUdj74n5FA5JF5ROaybG8GQNtvG1
a0XQ+jzdsugbCIYQ/u2vFuWZAnsU1p+/RuFjj9a2gS1ABflwqGmr66A/bVS/RrS6Wt8utOvKskpi
w2LmiFTUks0m/UNb1bJNezfNMPina+5aUXzioTNmYpVRktVeHGIVXnIMHTWNYjwfSFZUkq5zjE8E
SQPfIA9FVcp20vrUJB9D4/Zsh1ryBOCwkG05FOcVxECUI0vaADBCot8yKa8oStD9Q7KJt5o8K1Wt
d+BNMQmq1LYmYgUGRuJpdB+iPYygFC6hPsfvhNTPt90P9yCRXGw/Cyb7CmDVfYDSTevUyMfjTYWK
A2FsrKNeC0g9KpArk0u8kmFe2IashpCVqKXPj+CW1CMWn44GgmlB1ofKF/iwy/C6D68WMlfsCXsg
25Z22F0OyGyLMjUXC3BXe/ZpvI/lPAr+jxGW8C9LfkAMHO9Xz6LCXYu4Z/0mLlTzPiBBICyRniYL
2M7dCfIl2hJcIEM6prVwVJdFQ1HyCvm8T5BdRkUZ7Wxk68Awq8xbA2+PPsaa/hkZcKXU+hnbuXMt
YfGed5f/VFzI+5fKmoDNV05MSQLQsLd6iUZ41sU7kE+VrtlhKoMFNsXNfmIY7TTCD2xeaOsLrjup
95pc/0e+LzwZQUkuJXaj3vK84locJXELayc/Fk8pO+KwU4Q2XFdKlp2eBzZwCz1ralJc3S01Rzrj
8xim19DlAsbHTq0UrpNvhlsOFkf+4VeeesRuHgrFLCkdK5MsnlWxt5vF68e3IktTZaQWZqDE+RKL
dHuZzqmm/lkWZt3A0pyy6mXg63R8WEz7Zg5U1Eh4ysY9TxHejPa5MYS2LcRUOCAn5z5bjmPL1iip
vays4s+3o5SjZ/02bHBhSSDQF17rfMGNEQa+a4TEt8a2hb4sruixHMa2HrA3cU/u7ojVBgxHwik4
/RPCbTkN5Fn5Jbk1i7VTqA4Ai+qdqLj9Ek+XfsihXnKfijj5eJlK6eMpmI7UPa1DQuWk/0f+yPB+
L2KX8oKMXJCEh+3qVXi2cIS8pwQ+Ngd7F52IvM+rW9VhhAy2nAFu84GXHozeky34AIHswTR5okbr
ON4viA7pTVXn2lgkK02tWhrCLWK6b3FgA267Zd1MhstoehnkKpmzyx46Z8A0bE40xL/gFjXzI6vw
3gbEF8WR6v0GbRNp78aB2EaIWR0u+RQsMq4VLyfg/SeiXQJ9dRtEePWHKslA7B6HfO1d8S9AoNPT
Fiq9HmRU6+0xFO+64pwreiqTp4hv0ufybQC4qdnztOCGpAORubVjFbecuPWrzo4a7klEuUSaFwjv
aO081imRddXCQ97YbGEmQ8tAmCkLvuqhKthU525GmAlWJNRFmhraPDXt/YtlwBD6QO6xyuHPc11L
s5N2P8xUwTOg2RCxygZ+un1Sr5NxesuAp/ioJ9CdcN/RGolckJW2HsD8Ed8vxodDHv9KmjaZg2W/
QhCM8Ywy+DVl0WwjH9vBpOGmnFt9P/I49GdD/Boc1XhzP7s7qoIiAE6/GFZ12EnmwzhMlP6bR4qb
Q8iJHU5g1kVffCPwLjM2RJnx+BPO0EsJJcOz78COhE4pwCXu6Jp7mogBGmLZUERz63ztx+H36zNd
JsEEnr+PofzieITtKBDhjn4EB6iQigW6TRVHb0hSQcWmMwIVAVFsQn6CBcWpaxhL5vPGoCL8MzBi
OaXKYAAXU6pyVFZxNOBWixob7zfkPeQ/YU6TVPMq2onvp/mbg788SG0A7Taeizk1LfbkKvpFVUvL
I76FD9T/JnhLSaUbzs2SQ7F+/1H3yKAnLHrT8ppq9f2KgHd5UVL9AV4cOwNrIyzQTTU55/5EkeXR
CNjTSKYZ+XdjGiDb/3387cKJlKnhcd53pbF1hcC+ijbRgq5Ap81I+92Psi+AJJkjXFCw8vtZEnF7
j0zr+wVVK+a33z+AxFucWuiWTCEpPd8M3OLRvE/27j3MW1QC086vzckEzwru4hOWKe89cYyi4qeL
0lwnY7hOwn80CBNogiEENiPM8xLgeX07ZuJEUSD4dLJNlkXW4evi7sIoc8tjl0ig0tZ99Voxw0x1
u0Andz0p1FRxIWyLH3uS239NRVZLlXjGXO0R1aphj8v3OYuevPcVr6WLuzcJnNG4dTc+FWRKx/3h
vksBBgGddE79jx3JZ8MgCgR9rciBd4L+mzXcQfHSNNWlKt5wFGdpIsD57ggKVbClt2hCE9RDujr/
LPVrM8ExM2bSXscHfKYIBWlburJ7WLMU9Vk9ITsTjko44isNl9h1+C/Y3QcLsSEikL2vhdPuNv++
xxd9hKD+RSQlt6aaczxn2wjyYoHq1zLnid2Grqwq9lp57KAKx0LTpmvv2T2SwD3jyqqqXmI0PkhS
lGGOPZewZ8IuNOAf+k9PFAhuUB8OE+Xul41Fft0LXbBiC9t8Qv/QqRIVyY2e5D9JgHEjSkDMvn3b
KbBEiqPKbkIxXlyituN0fHfcKT4Rw9rSXP/naYDNOjpKW7Pzi29cbI9IcumcPMhaOqdFq4GOEBkU
5zoRAvxHHO0EbfO8/vBedkpg7QLOv4RWC3Cyldo0ZlOUTkRvS7ZQcjsZYIGB4PddYtAbYtirSnso
Jqwpzm3ojq/JK6I7JkfYg552QNNHtvZQJ6hWP4s4WU3GU/EFN9wThi7o3vtnSNs8Eh/yJxwNv0Z9
Om+/MZn9ql5AQZ9QR8fIGnOdvqEKK0GRoQa2cImkzSdEniOFeM3L9kNAluJQm/l4Ap+hdD1+88id
ojZy70vrL2/DRQNgikxeBZq5XLQeV6QytEfOX7w8DxgeNMWYtoCv0829E4I06vg3SoZOVDPYjobP
jVsEUVaCz3AApOa14PER6LcdQTFLllWVAr3HQ29GFf9Lliz0v0uR9a4agyrMMjd3ttH8XPF7sAEu
61AydOflyiZAX0rNGP3qTbeisxn470Z6z5sh08XsVwE78SSpdCSyTstdJGfaqB4O7FVAUxVvDAB5
VZHxGa+EkBLoF0nQ3F/Ox3tcz6hH4FjcYCSke0Y7624R8Yv82jbmS0Upin8XPJfRbh5fb47C5amO
WDtUXaC9CvFK9TktIDIcstcn6FhE9TFXWBgRGsi9vsTSQQxyj4qm1y26sh8jU1G6G9wwE34Oh+pw
9Mgwe4BAvCKqs2gCJfPfbpi21iTg8v/+GhDofJe2eOggmLwdhb3OT8dSznTM/x2PiGjtkRDg/aQj
49y8v/VrhXkNzajZxzoI4wAz2sZWNAMCy8ERzfBghGJfUBCHsJdJX2uyawcByr3hdAqA8PzQW5dp
uZVJfBmEZo5oDnL5YSIXLt1Wak5Lv4awG83cCafbgz68VmHO+XKP1U8zmerFdr8ke3RAJ9t0poPI
wDqntTmeHg1a5WAvorAHBVpbhRQGX+qOxoNxGjUWFk/VQr4cXV0iuk5S99BlPWVqMd+wSnidcE7M
GrYhpPCZz8T6lCEzlZiclO00r6gABm0RksLV7X5bV+anHwnZ8XdL3VimUbzqT3h9o9Ub1KSEM8U6
jA4cN+BpfdaKR7suOqjVWtRzzbe8R5zWoLZpKa7LrKct8ggw35AQ/nuZVBRGtcA9HwJyVmV+FpgZ
uKuWqVGNcNhvMhC+AioPCTzRtzwe059/8pJLiqN7tpMhT5NDP7Wz2MXYn5B7BkuOWXs8YX4E2iLw
XYaRL5t8979GK6Z2g6l96CwSU/9WUqT871IPj8xiJhfQoSTtJVSftoM6a28pMuYkmZzEANI7ShpT
cQvGS4N6MlrXTKX/geydcW3vuHrwelIx/k0vJfMC5ojDRlPwIpZVVfrv1vvNpm+ewoei5ap/nFl2
OPxvS/ZKh3Wp3erZ9M//XIKJB+8g/nUDC0cYZXPMEwvFODM7HCVBuigDSGsvWJbDsL2cxzuh17np
4vRUTco7/wAGXQrW2V17dbsEIwnK0loPfI5JjxnzdvnHaK/A/i2AAwPVlf/LQQgRDrXCU7fDkt54
CMf/KdEGTDzRELwAtoWO7e3t95ZUMVZIR05JzLLpsBd5WHvsmsmUVH83/eGTMIMVv0fbyvCncgx8
UpOT/25le84LY82u6iTQtmuo7RM25On3G+W2YOgOIFuMg7wMQRnqTfcN3dr5vE+6Imvcg10VDchN
MLQJVc5ao39LxpnC2dAh72VVYcZdW5OU6/J35HUuyucQP+kBMwP/mIR5xlpC2Z1lv461wvKnW1ma
ABli8oE8hi/ahA9+46GUSL8TrNqJ9EYmTu1wNpmWTGRtTlb5q7suF7086hpIxRitfCKkmLZSLPIb
Gdlv3FOOshfEPtibWW+MjJCQNJjqJ9h5dIfkFsNH66iEFgpSUhAlfhGQvmI05t/W7qi4Tk5ei/Jh
p2vpszDx9VSJtl0uPPkKUY+pvsfj4mrIlEimNftZLEUYZK0uDDkGC4l5uZMZofXAT9guNIqnwhg9
BifYdLR0lySePNkFfkJAjVr7pLR2mZLW3sgGJI+rEPPnLvtV/Di/X3M3HbcMJjb3HIzhmRAqAjkf
FaxdEmFADBM9UHgQesqJ3qPRe5XWez03G06IYg/qrOQzpgpsv3KYDiSqIXFsRqLs+gBWtjUOBj+r
jCAyUVgQgQ1L9tonNW0Z0ua93C5ejxtudPcAmHjgHMYMDVIeEKyht+iIL8SVArj/MeyDj0oUO9i7
b0dQjKn7gZemavznIRjO/uX6P5rNy4K4ImubcOHnPUq9o4g6bp0AijQ7BuENukaMyWHJmf7ToBUq
Kcf89Wb15Ph/efDhPQ/xW1ZB/52hi8Lyp23cBRikEEgmFyOIHOSvzbaNnquks71num7u7esANCyI
jG0XlJRP4C9cgddIxu7UDR2E1GJPvbDl4DolJeM1R8OrEBgOpDDj1Xpr4wdx3jyoE97cFnw0a3Y+
kNR1dfUS8XpaQZggpnXqS8FeS88lR73Hcry0W+1F1y3IOLHEesneqhRfqKRNp+RhLzdY/9PKIg5T
kaZZ1/bgbha1qUTF/e2gZyA4h/r9zD1sNO8cDXC71vxk9JdOY9t0GcFyPci1lj6IxTqXkTE8YRGn
9RFuAgpE3wcBaN5yMgfzkUDHX5P8kKHyb5mEYQTbtM7vQi9TsNyvjB7UQyrpyFFKHFqKGmkL57rk
eJ2o3YVyxBfgumJKVMy+ktxDxnOvwUMCA1slAKn8B9GFSy06kTHXwJlGq1oe5G7IFmvgeDXE27Ok
Q+oOHynoD6d6kRS5R/wP6+xOgVie4xTKnutbkkAGCPZY5O+6Buh+dwwOSzM8Zg/6Xp1K95AhZQL2
T/wL3k/vJ3W+P05ooIAKo9XINOP4v5fILpbJdKdQtrWjihBUmmI0QIgSSRosuLgYE13bRf1Ct/EH
ZRtw1epPQVpTm2ZhdX2xqmc3utW2fhUOjT/+FoqkAv+G8YqQYqFNaMjrlXB0qwpVKrgIrA/H1FyH
L8AwOawVkjkkA/dTLrI5yYs/12PsCBGduJNx2dxgcsEY1o+V2mPp0CKdDT0RtF/Ff/iwxh5jSz23
3i9g/n1BZNpJQ+F0H4z6FgAgPg7LoyRde97sNw05V3renQRXpRyR9QSQ4wxEd7gOHYKx/4lK7qQI
l2ZvaBO1CQB5rvfOWe6GkCemP2PvHFYVY9FgFQEvWyvHhJCLFAH5Q6ykFUpxOqqURLjvpkQ4BXtg
MxnYWsc45jDUWIBDIGIx5oKaHYxCWKNlanTtQ0Xy20Jptgpf606RgQfcEAAadviVJL2RQCI95Gpj
ZHrEcy0PAdu8zITflzQv30kIfCRJwHVADGvmLiIlsLKqfNjHzdVBi1fl7s/Nqr1kAipImzztIYj8
LKY6VzEkRKUIBsbiCXeKuDq68sQmuVVn3TwRnwUe/G5i8Hkf2w8XkrSY28qIl6fy1wNpZ9pIWpTV
Eli3gF1NW2eoKT+I+6hnLSq1yiZNw1zoqOJx/yqVY0dUud5TDfcx1A33PMUp3jih6ASs4H1xzQGk
HyWzbUI7vMnHJrjndNZsW2O1vBl474yCFtdqsKFd+Is5k1HyS+D6kLJKg+43HIbf/He67xjdWcHX
OEN6wzi9M2VPB8R+q57f/KJ0MkZrilYkCmSzkSEBE5FiOgJvNuHL5ebVKRDE1nFrAOaHEkCokOLG
viPivsVYGXH9U9c6lJdWiF4SyqJz5E47HcCKm+GJRm/czOaHuOeQvU2zCEJ72oqLrlpK8g8IW5RO
L2Lvm7HoTr0+0Pl2mCOLo/GMhtEFfJ9qvU1P1C18bcap+i+s2I/QA3+je50koKWE6sWqau4WBRon
NztgN5Qf0n+TDqCLymckdWqBJHHYrW7cwtzACcMO1uQdKg92i5/W8W3ZgUAS6bnVO8uB7hp1OIUs
1OKHu06Eg92BQs8ShiCWNhUx7MP8c9lp/zKNmAwb6kLrwHIwNgDGVqcRsFQpKy9opZmqnh40O/IV
toyk9QPKangkRotsChOCBZSTQZ7DiUBnqYR5pWHSiaKeslbjNm8pTLmMuOpOx71Kv3r5I3JcdcSX
D/to+TPedbiquon/t+b06oD7ymd6b74zwBY9AoKaxlicHgr1SEGLxMS3I4WxIxU28xdgEp1Eqz3H
ZdKBbIdF5gMhDBYswNNzg0an9SwvQh4oZABqdb/80iFJUjEPMc8PuIvH1cEbQ1iLICACsMjl0KMV
qOaLLxnZ0B7IYMR7fDuEbt3ECsSFMX1yw6y6aj9unm8Ez9r/z5txLb5LZVV5xhdv8kRJo0nRC+lY
135A3KHm8nfKytTVZU5MF/yZl+nBwC986WgZOer+a0EK+C6eDfL+rhAWSeWG6fXj5kWSsIFSPglz
VDuxUCFiZnwitAYOUX8mZb8sohdFGUJzDE6JxopOdTPqIy/O2TgH5rTKjod5QySxGUbrcUXvKFZc
jX5fHYupwGo+z5dcUUVq2hj6PL/ZKclIdk5Li+cv/t6qURVteNxWtqp2dUI6aE+JvoX8ybBKVqTd
S2ADL5TGOTzOf/QXvoaQkhN49W65AZd2PRYNMkP+u5qGoDWmI+773L/QXIcdPPB+VKMblp97VzF5
I0K7vNN2DcKiChznn9GMyVbvtocjaEV0Id0CQ947/hk5EFqk2LJj6QfDf+NNCveIVrukoz3xVg5W
Ce2nBuk5WGxdT5E8lOrjbCSilRQAJno0sIKjR7yxLZQKPweTc5CaUyjNnA3Kx4mDJdMEoQiLXCfn
0797aA1MP49QKdytWr8h+fG+3Sxrn13h0Jwm+x1sMZZjO9kLQXNM0MIIjH6ZjiNh7D9Ua/pGrf5Y
ydlbHogUwrrxi0wkQFzCMekA6HXUIhCWUYEeRLMfS4My+Lf+2QqPqC5RipNIAGsErXgaXabTkQMW
ia3tvank4OcESDvExyZg7ZAYK1p2JZXxO4bhIXLkbbiAsphdbiWMx+aIHD2ogtEq0vhCeVYUBclt
XiqJIb/H9l4IAYxkKJ/BSPKdy1G/+wHFOe0V17+bmSsWtEPb8iNSsrYVvQ4VaJRCAmggtRUyyq5n
z65aGTXI3GBaVw9xhw0KzDmD4QqkbNyoeH4E1NRT4fco/MzchtOEwpzwz0CpUig9FQ2ru8ZxISZH
0EjD53c5SsgF7BER+hebqpRypRunsfvSUSImBEAHYVDCeF/eHuHFjME4t+geGRxDp6eHKKfuBgXH
PxQLcN5nvM1nXhkZ3XDsXwx7wtyNF2MQSMbBqNUNmN0L7P0fbP+2doGgWNEpixq5I3axYvIM5WJ0
ef1Yx3VdtM1PK4697SvDDEp8fPRO+y9TFh/MI4nqtd5L+/DpM9dd6jfV2e60OezCAoWwiD04uVUQ
l83cd5LQdxrph9NB2RmCZ/E1AAJDP05wOIXq3S0njj8gCKYiHA1wfdi4G3qnuH9aoLGvXq2mKMhY
SUF07PpnC6yIUz54BG1B2RTYwohTe/vxRNjnQKbsk2Q9xQY93OsK4CW6ggQirpN+Nx9gqKJZFpIW
4KerEAIaDv0dEb45smB3qgFaSgki5Pf7PDoooQTb9WCB4GO7YjEd+AfjQ8F3II3OTsj0rIesUdJT
/oVjc7KxlBDxkiVDnK8viaNOpuPk54Dbpt1zFJFagn8wMOJy07i9+rSZMOByLuAn71leDrcgNxhN
93TsHdSqOnJKZvg9fnPXoKHDCKBclefw7FFPX8gvwv6VK5Ty5BJIqeqCosVO/FH/+ocy+uWlNIKJ
WB79Q0w+Z7hDAPxQe2TiNrddUpa7k1OZXDUFieVm2T+ThCw0nVAUd/pGCRf883zNq1E2LOJdjWyE
ArLk+OzvcOXMdyScTivoNMjCIxN/D7NH3jPZI5im4qME8VazoDWaaRaaVbsC3xk7mvespqJtUmT+
KTK8cL8T0M1yeZ9m5PKHvzsv4U978pmWGeOnJBEfA4UEpNSmOhH4ScVq9nu2/nm49Gx1JMCBKmRp
Pg7rHFb0EO+ZCxnL5howtjj31mkiLR5AeWZowm4+t7ZwA04BFoji0yjD1sgh2STZIEAL9vsCMcnd
EpLin0X38QFp6CkRMaGZBrEYHgLuvdNI1bLTbadoupeWXjoJdgjP88LeahZ6dHxA3C/6aUAgGL8W
BHzKMSjsR1wwEWFNU7gTp009kKf34qJINbXhS7NA5blffwdSDRdgiaSHAXXCpzigTfRgoWBumqFF
L+W/dHrcgsOeracZyQ68xC1qqC3U9W3ByY+qw9np9bJ+uiVyymX56ca7Zu/0Cfz3PH7KiCmqPac2
hab6lWPMhf8Z+sP15HqUf/2WoZGz2M+IIlX8CkZ0JQuDiDdyzu4oxUCaYOp1qTaEhySs1CK3wAJf
RNHEZCe6IetRdhW8T6lp/EerfxbqFl7Jw1DxUAd8r4DYWBcPS9hJWioYyH+yEsIAwx71XLmVXOoY
H5Id+mjq6o1lSj5lJ1Q79L9DHZuIFhA9qMhcmmGhcO1ZLfJApescgGX54Q4j3qT7iB3FuC2yaX+/
sioGx1VQW+KSe2POl1hgTRbyT6y62qnaE8VExmcuUFIqaC96aBXFIMa5aXM7Y/ModnnULT0nJd99
7rHY3Z8O9nPYHIo3YftmnM6Vo2rAP7ZMb/gXlP6F+7mLRjM5LRAOjXqSHJ/JCl3KDJSwwIicc+60
WWbi9PPwlEw0Tgxvdv9g00AMiGN3V7YT8TVzVWqNK0Hq29sMVnah/2HOuh0tOwwqj9rF3tpvun6T
YZe99l1U21V+6gAhcJMEV3mIaMPAbe3SoTA322E9A0XC9zcMO5Myv+NsLZ5IK2zsCUceNBZfBlsz
F0rJ8qrZA7Evg0XeCDlo8ebxjEHKPwoJom0cuUn6G6WsCaO/bQv9JAxvbJDIA5YWjJebK5LW7AZx
7aBMe0JshRkyfPAjFNpLZ7+FK+e5t/tqwNlQaUixmrvsuCEhk2ZF8ulyNHfUTdDK2G1QQGiMz4A5
pZ1iLtIxIYW1QwkH1TEdNp0dZtrOvh7HMlpLr0qdcz1ieYbk54w70UKkpGMn30JkeljgLd+/K06c
S/fjejwKblna7ugO65iMRCkjOIeW2N85fkz/YGEFBVHLdqz/BGERi/hoiTpU+NFOjgk20EIfahDy
EQ4MzhgBt9baIPSf9aSzLZ9VjWw7417FvjbHVbuo5VIbdisNFCa6qgEeS4qfst4fqBUVgtWMHjIy
oA0AD5H6qbTyypX83c3/+BCxwdAtucVjdrZpK5HY6Drlf2fMvj4MCpJjDJBgQXhc0jAc3LzaDCAt
SrZJTjm5SH7bErdliTkEdm/G8wHcMrZoz+moPcesnujaUy2J+9NQNDTqhM1ApoWhjRywodreumFs
cRBroQZdtn4KTPSO8uEu3Bm/onLQ4jbbHp9qGoaq2jYw8bS9C+tqs0mVz3udSLZYumqQr3Lnk4Dc
eBUyyH13nO2kjrd4VCOqGf8rgjeIqDcrxnfMLfh3U5TnYWDX+VQwJts6jm9M4kk2Loq1TxAyqxZh
xhjdgkoPIyJ/1lMWqLv//EWTRdkCPl3dgHShgjMaJo3lx8m2bpwZ2X8rbaCbKvwMS9mdI/4+rsE7
6kIKPL6zF8fAwI2xw1d/LlFvWoxboDJG1O5kwgarGlyyqR1oabBw+otJW5OREndvtIWhqTi2BBlD
HZ1e6KCvCre66yzTEK0eFxQS3W7SVfrgtwhxiKMYeRnNO/Tu5an1o9HSOhP7qxewCgfk3GedbtUq
LZwvfUStTfMNZ/Z7sTBdEumLCIfkjXoXmVdJXNhnLoeDReinAOQ7XlnifLFJcyKxoTlwDWs6PM+O
CZhI6zV1OUtwXYRn6qxYJeWcr+S4GegPPMCbZDNcUfV+bGEc0clLrk/qqBuSMNBnzfy5bTfVVH/T
AUGQfdj/0J8KEdzQ0EWRw+fZTPQrgVATqUKdNmDoWYI2xKZDfqNeJMBUE/NRt1AoJdqfQolUe+fc
Jy5xpefVwwVbENCElZy6YAJAF+hFzv4Paa3SqxKoLokPkrtrjN4ODZVYS2Lz4YHrmp8g6hcIotCH
bdu30L0+ZGA/GPpob2wCPPvLiG2TOAGxpvQ3XH+rYwawh9NJ5WOaigEN/1K3Ij+q7ngd8UfyJWBr
0kudCXGxZVfEvDM7lJytRQTMW1vhDTtBWiX6ctcqsbo4IlRbkzH7ThVAR4l2GBa3wypC4Ie4swyW
BxjXIkSvEpJ8UmbSbcdCPesM9Z0ynZJEWjbSu+wYSFovz8HB79zHv33fLHNdxQkebxL9ZriZu8vY
E7kzMUmH8igL15aKBAYmEB2ittyjEPC0Steac2AI0v/0lImNbnMTUcaPy4LISSsn9jAX1YJj4zev
MSJW0nojMiqjQRAedNKy7IrpOPxkKkEKQLKPo3h4fOQyX5pGPdQ8SXbUDIpxfGZR0HChXHKuYL/Y
t1HY/2HYxyQMIk+5TKOTJQPsJI1AqKHUMPTCTTvwtdxXIRbGIKgqFQhv5n3lr7/3Y2p3lRNvDN8B
dgs72wvI+4QWFTeol8eM0zzvx2SeTzH8kSRr8PAe3d7MjgLHZVkyVCreCJ2F3yapngp6wqp7VNeK
Ff3WUZj/yNHjbcEiqKpOo5gomhSupB+bX0lq/Da122s7PKzovC/pB4dEpuiccYWgtvebKFRxeju2
9P9F0Zn3Chp/5iiYDABVPjP5pMLjHWujPeq5TzCBCCbN9dvettwde9gduzQWN//HxL0utMwa0+HZ
iJ/XCaeviEIJPXff6FEkgIARBqSDtvFvSNnSoedQUzXj67xP5ej9aLo/dti1idinGECJHcUGwstl
SPYOhllh7Z78SiPOJNmrHokxWGOz3tc6x0Iadaf9q3IvQbyJvODQ0aU25poI7ukzZJCmnrbkuvjn
ZUbBH9z28NLyJt5LNBqncNQGwcAMdqaRfA/MPhCqc++EhePzFZ3V0wg0hbNOATY9A/NhPcp48/ZL
vk+stWg1TZVZpsEOuyArrpzDzAatEvESNXBRW4ci51R5a/tdtMVMqaxa8JeXu6lWA3Qp+RVEUF8C
esRMQIDwK36LZCpmS9qG991DK/+x0HmPT8jxhuHD4UXlxByYfGYb29PyqE2h8bDpc+rdDbZcApGc
8kp1tnHxD0zblSyd0AfKPWcx4WcZlCa6vQB64lBwCtYR50zejSuBcslFtd0u6K8J4KUPskGdQP4y
4Gx9mkPU4hjrYGAY6IVxkztjHBMD2yG6zs9+p1fhK7TiHaLw4KwcpomucGjWIAi0E8VkirSMMBYu
NzgIBAVkDyF6X7Zld19A6ORZqefdnTz9RTHNsroLVUW5+zKVxPC8+9EU8z0nFZIUKmDhF0gGTmK8
PCB02sIk5CsOVwTfzRyTG0GnWUpc3l0Bz6YaxuR1n9mhBYWSv0vbrXNcuTZ58jlWlzjQp/SgbqE9
qftZ7Og66lnSEiK/s4k5pUeWakvpMwa2Wn3QXDyr6TCfm6vHM/WNtV6aVBUR6+rG8Rxwffs3tZIG
giVCtqQEZXH26y2CHkYp1mWsSrjYoZrBaX0xQNk3HZtX+U1tugqiampcVdsxc1mySoo3P2iARVCC
Je+Atj4WEBkEcUgsz+zPx8gqx4f4D7wBD1fliAn2N42e/Rj1aC1iZ2iLvpw8DHryZ6UEzPZUY6XA
gBMDX7EiqGx3FowBlQT+BtanFU06g8YTzfdSNEUbqKry5F3yC6KpU9KaGFk5ssTIpWfITtZIdy91
iU9SvXCvFic8qqihPnml2AnJSXRJXGjk0uLtezvctwJd8MM2WA2Zeh60Il1/5PRCxDNj7qELEVJh
xZ9jTh9POaQoE/KPR2NqhqNnK+0Gep9ivQ6bYZm0WYoZmbI3L/R7AO3iXNvZAxUci/VJwqIt/xvI
4BLbBsukEU8wNSZZIbZcGzprh8LvbZ8cXCwiub7ZVo6CmEoByd1X8iM8z97YnJ+OOpVg9vIBjC4F
BRWSN85rjQs3AvCx/hyMIFheSkXIMS+L+7+kkWTZ2zS8pRgbemM2jMw4cj+S3MiKgJZUIgeLrl+i
07tq2X5H4b3syHUvEjtVri/9sbOBD9XIgYQB+4cUMGckCTDCmp+eyMDRAnecW9Fpcm4oiB8fPDDP
TN5Y9rvHyXvg7wyPl5gRSE7tl95QWY4Lu5elhkAhtvekSMLQ0Lyk3HLFFS3+ndT+W2c3TQu2MLgY
q+OMkIQSQwK7RauFn+DXSdEG7zVbKgWR81hNpkdX8TltW0TMmAcHHTSirbWrH5NpEEvKDPgoG9P0
oYi4TAEmDkJACCsEvZcE3mPS+MqhaTMQJzWgO6xxfja4pov62sR4FIowCHF08AqGl5UNzGpUx/I6
idAeGcQeEuPKwf+pv0ew3PWk0lOt/DEaBnMf0HqQXlVWUscJNnfPLnuJTjfB1XDW3xHZ3h1ST+Dq
11salu8LDuUul5oPJIkUFqVu0g6Fjjpoj4PdAYacFRG1wk54hK1QAlZ56K9dB3ZEiYdRRuXC8+hr
CYV83rjioz3Sl6zBZOm6O5y2zsQHk2Rzz+Ot1IxZnxaqX+9rzLw+bjMuuBZ1fd5p9BGPtwApMZv8
LJZwGzRiWI+LQzN4yPsUO+9iWp6kG0vbVC+2d0RhCiKLkp/XCTlRloqPZXJ1DyfEJzujPqBnVlA3
BRlycbsmE79F9oNwx1qgknrFSoGd3y30Xn1JtcyyfSPktzAQC0kM7RxnOP0vJ3Yabh+pMKusklkN
LQZA6hEhOr9gnS+P65bQtBZDbr8BjBnDRz1jY57dLJx1QgoS9uJiQm9PeWZm4XXqbCuwhfPtHaMO
qjtXuBXMkDrSusnBJVlpGrbY9b9eXcnvL8x634Ve0dJsney2Jnpk2NR022ZkUHnRH9uvjRBNGVtb
W8ONJ10K6vBeJf0qwXyMNfxwYOCjdMTHTlYV6P0iu5nJ+WFeQQAEbiwneEYoBE+H7CGahrV/ZbgP
BmThRqaCHq2inIvUkOulkPUgHgk+oRIiFEeREgqfYy7E0BMu5HKzsVzAhYcm1GY04FmvLdKc99cN
IW3jqsgBQqgjgfvWuZw8OiRHddR1VeK5FXhZIfjvrDdOV2QUa4sCK2Rv4JjUJ0EalqZruiL1pqnf
25G3Yrf84CmwYvSw2nSFbIgRs59CtkPKJiVqrjXQUZwRKbzrwZ0CkyORd2H6UrdHRGOh44BoeR5M
TcOWjW173QsTFFeRjqgfFN+yHVfSP/yVYc08gUMD/puan5Pt54xbHqg27PIkQiiMeO6f1bu3T1Yw
63oQV5YK+yBdPuoejUtNC+fqxoMPmuBG0RwLx4YxxrsdKLSi1++XG9YN6mKlDQ/9sI+rwmHLp5cT
bSnyHi+vhWhvBWu0sIKQB+TwLWmpUvHWBf3n/kHcBfKwm9aK/pB86fNqbeEnkH5KnQFof2wkpfkG
H6x0gRThXiWc/JXtNgmKx+gaVW6X3Ggpdnu73KzyQUnTK9pcm05jF82tk9CuOj8rItbUodq65uSX
kqSog5a6iYAr+NNfzEIZgteVsXJ2qSvxo2c/XjhFEj6AutVXzSry1haJ0ePSCP7TLqel6g4FSXZW
sZPF5ZzMzbG8qe1FYvnJj736GW+YG7Vca82tKO1PyJ2hSH40NdIZMSLDeG5V2zTYF95e70gJLsA4
fNwjA/ZZjg8XkfslOMidWdycmEDkNsW1nwjKZXCgKQY1BbyffqbJ0mtrqAifUCssl0VYKOh2xGhw
tyS3xy8Lf7U9eNnin64Oxl53CLRvftYutPqToRZFpRcDnmokzNtLwWYX6Q/OMk+OtW156UiWtOqm
DmGTIqZjB28EP5Qbz5+dkW3gjoO1Wk1o+JuIrPMeTiNj6W3GyN7MUF2mmRg0dUGUH8DqsHRBjs0b
rm1bwgbS62rju8Cgd/nrWrX714SEb2hADE8rywDeAbeIubBjHHVMhxF9rUglgWWxUzmJyfW6Mxg2
IqrqZEZTHtcHQTHEy2VqYUx0HsmwRssFyYXB2F3J1g/kU0YSf7hj6z82vIeE0CmSfysNxTH3ZlD7
LURspo9ObikYShAHgm6RL9uSnw37EA8WKBiGKIGtovaYdGPVNZs6+YDl6GS7DERV3rDOJcOlONGj
DsgpgT9ux5QRAYgWbzyKJVvI1Pg/j1zEBPklalpjm8qoG5c0ZP1Uoy2n72gOPEYdI8W+jcvpCuHI
WxaasDOZsR0F3AY6wWHum4Kod7QKAO7IiTVqudMFDjgdqIkZZt1aIs7S8Cr+kA+hLjUXHb28t9eF
asEP7jgdZXKdVlzSWuIiOb+wFZ2VzYxcHzY1iyy3v3vRISpxHlXjedlOl/MJqG/+vrYXjgeGpn/7
BR11+DLmXoP5SlVD8CeViSW68We5PN5qpaZa/d6G9zdeUkMEcqCkW2xRWref1ZRhpxUs4oUjJmPF
Pv+FFQ3WkBFGO9DP0mSwVdlnKo9wSCiGuwmh8WDqceZobTZyksVwPwQB0vlS95lTTjRdbgUVJcmM
MZpR/tMJt+Qt8hspKwTDeWhATNdNA03uhFumC/kkwIrUTbixOhQMtYwHjI6NjLgo/J4+Sscm7lYz
nz2TAzHXiTKNkGLauRDTrqWbH8DU+5zgx/IhaYg+0nlkSYpxXV+rXgUmn22sKpXnPu3T74WEhxBz
IGIWN6PvwR8rPOL9JI8bFcKEZap6Lii5tXxhoiqGrIhoAiUQsB6g752fW+qXnklqqbTpMhTM3kea
UUy6xV/5hNjG9+AD+ZnZJT6Lv1/dgrE6elNdXSeLpU93Xb7frIz5FM0+FwFNLR7SmJqQeGGp6WRl
8YBJVS9FVjdKsEWc07RIfsM9iilbdVbA/+5g4HCs6mDhsG+hCeMbnXERAcwnE4XEGynOEjHtKnPz
cJ1iB7q7yTU3nyrvv5OBusNaxzulO7t3xcBz/EPyQGaHJ4UNUdPnBs89p+E4IZUF02CtyQoGL9iT
XTXqItQlDxD4zFD13utFBk6FEhHbANofHXM8hfC2S+xSvtCHUtsaXXVtAXV48vqBxUdNK8DCcgMa
lmkEFzqnsEFEIqu/Uk7uKnjo8OPHA7GziG65o/oP48fQ+YTF8bCYhXfACZHH+Xd4vsgHthueWPhO
+B9vNuBzxNzUwaL68LfL20QRCPw+UG9q3B/3qzzzn353LBKu/BV5YQ8bnM4SOhIwiugoylaJgmPI
kpuA24f4ymDCbD272I5tuGwawhGmKMqFXk7UN4wkw5duNLUmo5jBsdi6fYIu6GFP+7Ndewy4IGyw
2HwOy1U4HBAckzp8KosdneNs5BC4fhDV/uxwpmBEEuZcOg1f4jATTYrfvCrHT6NzrEPr/eYj/b8s
k15iyX9eKjCBDbxP1T2OOkhlt5bwVdAm9X3SL7HzAT0U0Wx5sFDM7R6PdycDwiOfGrmLtXo/1yJR
wtu7lnfa2rzqn3SeefHItUCZ8RnnUqPANsKbXB6VXnnREGmuroJRdCcNzWYER9o1jwJGIXxRmXvE
B5RsBD9cOwrUJ8o64Wrc/j5qgC9Ii/1M9RP9fd7rMa1ChxA63Z77FlKXo+ataMsc+bYE+C77FLOO
IrcnnDPS7BQMHi7w8LX03SjE7rI7IVi59cI2hj2JLzMrshFzsIDfvFi/YPiT7oExI+yXXFavDMYK
aGKA7QTAaSWNEDS5QAMdBj+nU/uYXPxdZsBI7oiHOrPT5gcT969yHrKf8PAhhONpzuRTNZzXARvT
hQMBzlpv8aEw84G0xotZEsMwChrWh6NyeB8TamrJ60cLXZzpIlt+iplpmuh6k9Kki5YhCBeSHfKN
gc3ICZaNRTn3fTuQ3/lDElTVqZVHmelh/p8g1J9fhlr/H9EiVFS6aDmt1ilSRh/yHKOJzGhKjDos
jOyEyPVmR6tvGpUzPShGa3PE2t8db0Nq53tuGxP0RQruzExG2sELH8CdOF44XcJdExiT1HEkwS/4
jToLTlXT4PGmQ+XCMQcfsIFxv9MqCUI+tAgcH9anhFgDILK+e1OtVX34Njn6f/AM/kWLnuYBD+tO
llTu+sGmlVGK4idHVlNOB69EetKUjqK52EaXKps26yRT8ZKGEpcTIYPAXXTLB9O6XaOSaPu/zeWI
cMUszYde+dstj0hbqWhEg2movZNyQv94gt9ozldb2n5azz9GllkpeD90G8lvEx9XsrHquAcsgZN6
zoqWA69GX3QyfQaTjx3ihLyFjb6Pa5fdAgM0HwKv6Nc2sWrz3q5WFLb1xDLG55MGz+2MWNV+8uv1
Gp5efYrMPPq032cp4aE0mMeEbbf+Zr/KJMvEN91kykW1XcN8MquCGkI/OaDB4nxVFTmxYMAJLL+c
DiFLi+Gy9eEP6MlWvDTPvQEhFoZTJh+tE6nQXqElsuiUsymc3RcEW7cEihXgromb7hy0hQNN4Cxb
dNSkXlQduhdS4czPPfNtppLVaiyAA83t4b2Qz95q3QzmkiZCw0PeSmOQ7Pj2BdwEsNtXe8fmj8Dj
/9eYHMdKDy5+q5s/HAgI0QfIyeeZCojAbgOSlUPX/a52tqdELujhJUylstJ/AKJIukjmL6DF1EBX
0nPC1oT/DLqA83j6eKiHt/CAdwDwnnmmiJjmop2RNKhmMSw8OQWwGhlKdhAGD88pCUDSvVG6ZzTa
KtfjVmh/BBsCajZv6lIHVSpM9EQHOeJYGyM05B1rfkDJlGPUTJid80/BaZqdbmG5pa2Xkd2s/d0a
LM4DpNJsDdh3jFdRD98ifOhKLLdGq1AQoBk8VNU1is+GHuYDRT5eFqeGgRYukQwlI3f0fSONANp9
wcWuuOmm7OEyRjh1Uq32w7i+U3SA15c2d9bhXEgtUUn1FdIgvB8U9o9xvctG+Gnd2bBDInNCEbXw
5oHLXcFlWcrr+ecz+DDszKwMKu59snPGO2Mi/t+zyTknQ5BPHLzbM6pBvPNjuO0I7M5rDIvHfKvo
oqWC/IE2RjsCYBWB8Fjf5n2Y7RgX7wgHt4jRJvlUPylCMhaCrncdn+DwPEnttuuDDNTVGq0gPkQX
1z46kE6fnP/qOniGm2VdJBVp0V6zHlhB1nOWuM7nheEKfx87sjvlQIW24aGXyAgIZX9VgoAXbpWm
vU3FvD3msLbDoMcVsC8vh+Pz6LdMfWSou2VrSZJUzZy60ykQBJhfDw6QcJh6OSo143LKNUq0URU1
+g1rztlY8EI6VmYhVN62biuSdcxYhIg2rL8DmxRHY15BleZZZsh3Pea8CN++huLgN4uGPBbEWhKX
xbQ+UYHjMtwvlveN0fFqB0nnet/5DkmeX1IflzwZknMMIQJ4Jx7U69PMo6b8CyJjCZoTCLoZZDDG
LDa3Iq2JJsQ87VAikwCWLADA8RkPpCDSxzlFo0BS13t2Inp+8Ojz+SdWgL+h7rit86PNKt2PVO/5
gCtYtbcnIdXmJag5fCtMNelZn8nam6jsIgn+lkysz+NcpvbFkW2o3kY6K4R9kNbBvi1ANTN2H9HQ
moMvZA5wtOBMgC9DEoBSd/7G9CmEIO5EezQ4Htgc2qN3v06ZTKZ4llkA3XNjBWZXEx19ZP7THCRp
/OPXg49Dht2nmeLUDH0jdNJQYrjr7rZ8MJlvB4GRPx0eAbfExipCbInra6WECie62dnKvUydMY1u
0alv43+ssLWl0RKLgCjLyYmm+oJdve873Kp7BFBsuIbYKqBmcMmUN6iwJFAJQbwFzxatGDBLpFzE
4wKGgPvYUkFKLsU6lx2Nhha+PXHLVgjhTwGkFOmpARpvcOjSpxTHOMC9edPmId/3NgfMfiawnrms
Zha9GV6tauzO83EjdtSCsu2bV5Y0q7sE55SeaN2TWLNzysheLRYHtyqBIwvk/zpw26wA06F2fLBj
IhdZ58b7VKoMSfvE/ys0UgzDSvIIcJi8kGD3j+0PEeF1hz/CW5An3bpCkyiw1On4mRGpHalpGglO
Vkl6mTdnXDK65CFLHSKgdZM7w3yxZKNYRnTDma/hsDW1xKAa1W3AjDhRKZU3oQ/uWYFhAlDnc1rF
ryRuWGyLJ8Abzwqf71CDz3JbgXp+uXi1khXwN8AaI0AktilCL2+ohudr0jL9chcZZ2HLDaWNj9uh
x8REi0Rba3pCGUUeiwc+UYTD8gRHkUijkSHn9icrx3KiXA57uPcRtg5DL/nysHqccrxwaLgPrATP
0jiu0NnPGQqISPUdLYAyNpnCC+b1HFscYvK9n2VqEJRjpkIiJyTwPQ28s2HmX+Jd0ctZXr6wgrGe
eAZ3MIdRc3R/cHYUTgT3UXsM6bRNraDC7zm6QrxnJOvLgThzn3uQ61D2/FYTJ7n+oOzi80U4l/Xa
HJlWmJtrjOGoQqMZ+O9BLYsPkg0iftqTUESBG/jsX2zmex2qaRwPEzoUF9/QAcIKg2thDLb+7L7b
85KPxIJpo9Oxm4aiAW9lPv0EGT/PwKWatqTyDBcDt60NcYqDR2x9fKP0JgQ5xbARRFflgCEiYJcJ
HheY2eZiFYBgU9AjJr8roB7m+W2MDIwlR3OGZ6cvUa2crwe3J6y1ScbzNhpH0fnvprmD+wnn8NIw
78o1Ybcp9IQHzj+DKuxStdY8SQnoxpXLJ56f9L5lIqgVDN+F2sXd/0/1zMqHVvLyOz/4rgPczj0f
vueMYdGwA5f3ALHdmlGFXIGwh76pvezWvrOlaRIE6mTsXBSIELuWvdPvT+PtAgA1RK2G1oxrUijR
EledFY7AYlLE3OVgLLoYFbYgNYqLkanyTHlXvHefn/RBOW2+mAMUSMGKAZfgBZwSnPGBJP09j86Y
lGOzCUbqrIh8snocSo/TZEcid1FgikN9PX95MbzQA4lV7fF5O2Yrdofi3UuFx2uFn/p4HG4+jmd4
5TdHT76vCq65I/caL/aUN05vuhgXMIyUAOqM55zk3FeQr5dFvNga8Et1FgJFxByt9DneCrkaWWY1
8luFrMYKylRU25h5GmD4hYWwEZPvmFJN170r4/mjB5lM8/CnuuJAbplv391TnKdjfkX6ZClH4B3l
D8jf+TaeXuKmFedvOXqIP9FwqZg7JG2HVdTs8GqlNc3SOcCTGqgS55i1MK0c79N3SAZKeP13XZeq
ShWjU2/uATq4OOCI5quvFnwp6Ru3XaFnyL6lyvfB8p5n2O1g0beiAr4ph1LGKRAf/qoNh74dDIVM
2kXFr9jKxH9PLa+Wywd91FRS18CSUcEMsXDBkyaOXtpgPOieoBJwAPYXvHPJ6A7hBEl3/2UwgOJM
dqQOnCrEbDnEjeXzAon2mPBPiMh3N14TF19aFvRPphfKthO8DTxgatFCR14Hn05cRIJ4wddI/9HS
3MczAaGsWHqNEY+Y+C0BwjeTh+qdlbXJW/dAQEKjr1oBf3qneEry7IpC96ERc1hZBPb+bLvOzhAC
8iLM4dowHzlOJSJGJQrYO25fiiR62pcWUVl7tlFw0uR7F9dOUBZrJU1nf9zw/rd6azulXtoTul88
E8+puCrqj9M/QDJqvO/gFeddvKxAlkD7+vQOQpgDZMQw+OtHWP6PSIeZ2b5mtWezlOOMW4p94FUV
4dL56IKcdUftueFMZXL0uU9BYavNaC3hOTW+L55akPqv0nOAvv45UhubVmm+/S/0Y+IlrTT4huzD
rzxIvS2FRlO0Q7s+VG5paIK6eHHfwwhQm55vfxtctJAvvPsIX81y5n5SY60CJK/rfHkbdC0HXVRB
uui3KOT3FJPvix6hE+N3H9RArxMqtOuS14Afv6zDFzgR0yvONqjlRgxRyZl8hFqASXnRZWdSL0h4
xhH7JzIZvw+gu+leVr0Rt7DI9fr84aLP6/49ZPUUHMHvgcWILl/A6mDbRkrIf3YjmRQOSJxVfKJi
T9j/znrtjkM+D5+0rDnBk74TA5uEk8Pqp/RIbCOoxU5F1AEem4qFMRc56RjhnAW+31M4kgRBnr93
jmRANgV4iuLBKIhn7F4YRLidUwT60N3uPgUoIAsobWW7TdnsoH0Q4UJGa0d37nfyQehhmQbnz6cZ
MhYdEBdzB34r//LueIosKMIlGKJ3Hr6uS+s8HE2tBuQWBNEOW6pSIo3dMZOb0RkQRVCGx9j+PIlE
qsF9TC3alCVwiTG8kWG998pzdvof8iiNRC6YcAw/iHkxL7voUXx5Ef6k3P8yJzglHzcdgQRM2lnq
K1NAtT6yT+DxdVy7y9Y7n6SeeRaaOhfFhbrGfN+5fZTDLE2eZuDDmRtQRy/AsXH0ZNiPnLhtyiFy
QdhLCy0W2+5Jqrw9hUUyigDiIzH2K34IAKGlZEqDUSc0/BNmxcZ7ZgqFq5WzxdI1T4KT8IDzHeJN
YHWmXHyq4Ttu1V5P6q8HwJM+ElfbYtZW51VB4uypBVEVFhF6MJkHt5+rp/70t0x5H0VdyPhAx88H
KoLEm4xKUipnZMBy2tsaSjgBVchoKtyYuDoV5QJU9zM9CubqqcuQ7wABJuw1ZGWRAE58oKPH8m/g
lmqjufKcz9tg9ASofICqOpjrqzOqvOb9T+wDnwc/R+UO25NwM6XAkUcInNTnbV3+6wBifp05jYxi
TdhV3OexsWUesiYGd2DAzJiPnKV9VmTTbipOGlME4qWyCiBFfdrZ1bv9IGrMiIbLUQb8e/vVmaE8
bN8eGi3LAjsSQUjRc6pday/d7jAHFqNNIM8gFGfhB58vhpzD271NzpaFn98Ce1eEdDtFd1O7BNGP
vE9+rz92JqYQEQqn2837X8DjOfTyBo7s/rs/xIip243p7zjvoWWeWOURew+e3K1fVda2Wddhn5Lz
LuVNrhkCeso5iFxytMsQOOHAoKSPdsn/XM8VrCi5DATcwzvhwG7bDIWmiUCc/Vk9n28R9iMrHT0R
mLKDU7h/zxnx5tAqdV8X6oGUcaSWUgiyk2lA9/xCejce4QfRA+u7lzxkSfNmZ8ScMncEmGGKhf0/
jFE4q4OF/9cZJGt+bPeCwoExkvLhVRkGzUaxnWtVlENnRtXDH9xgqN7M+eqYDH937TleRwXGxun1
0D10sB8VhWWqG/mNWszUXyDg4lliOGgvWOdsGcAPASSK+EkXsPFs11+RmtNoWWhPtHD9qAUO2nLF
vEKgfKHdK1JbAt0TAVNxUQYq59bsi/ZLsCihEGkDpuJCHhrbVGP6mREVWCwjn1MWnk20EGgMxTYn
o07wZVjNqnZrsPD8qvGUpNFNl2W1jSL7ahDDY5BNuOCz4R1LjCYMGl0ZNIULHfc7tYNyQnWulEMB
TMc9q2/kq3GumEhDRdTsOiPcYTNSi1NRn7yDNq5RIhMm2j+BGrEsdY1KewivBjbUFaQpYtbVlUbr
pQ8wEBfqWoHp7SikqVJmGK7HRZuUGTu1x17V+5tDXoNeaYOOztIr00iPrXPheDnB2xOHdi+veh9I
dgyUlCIkXDSuyRZwDEo7jj9kkYknqHs1CIAiSSceyWR3py5QCcoSW7d2hO9GcggCDnhpYagGSGtS
pn6eech6Y92t1KzTQT3nYQL1qNRF2/9ggB4oog6Le0kLFbci6vJfeMLQDGHoXXlpGMsmAiohpMdx
Jh8mt7yLzwaMJy0vLGjum7kXXs1ahhrJUpVSIO+bnLugNNT9IaHnTb/BmUBWiXEZHI/uoVOuwrKU
zdTk8kZsohynAxdH5onnr9J2bEZ16IMdTfs/FmPhryiJExwPEl/joRhV6sEl3V6HnrbQTA3ljYFv
+bv94H2ID7m36K6zlAC2cz00D8grQAYJyzrah/gG05jAGBwMYjvzh3yUCwmrnfQQXjpQr/6mc4i6
3dK+CYdVnO09T5O/DaZ6gnKNWlQbYInrquS6YMJiJ/m6hkClrpBUY8yXfMfQOuOXok93MTM5ZgjJ
9ildYrcZoZsLqBfhhi43YK0ATOaMxHFh2FbtPFJ75jUUeB3ZZC12iGasdts9AH9moCms4Gk4JLO+
evaorpQhPIwrKGqsCMOQTSnB0LGgsWXOn1hRTOrLhols1CC4u8nYJkNh3lKvEKPT4sDLBp9inCB2
7XtUB3pqFz+rVrghQ0lRqFiAhdkfSytSYpcmkQdx82i0KRzoaX+3Hrzno1Q+GVuN5qc2K5lW32ss
6TZbNJkGch8tEgZHpb23NJAbn1fQaIy4VT8+lPel75qmJGF+tP/XgX9ZLQiWI/3ISmZfewHHsbJR
aAgWC09/SOTQxsMo4Vr8zUOL0OXjUXFEEYKrEacYRzyXmPAarsxdhQu5FVC8clfxfsvWYiNqc0TA
JK9shz/kaSY2v3zl+mJAzRoctG7j6v1sThu2w7cWBOBbBwNh4WUM86Mh274cKL8+kG7mUzs94UhD
DtVxaKkUabM95WwFDb6BRuzOHjSXWz3tmtKlp+TYQKpFkjESzZcpjKeq37R0G3t1vODfbmooJR93
5/aGIONjwH4DZVlAoh4UDoXqcgnilq9vIxwBsGe0M8/4PX7kc7kBu9PU+wpJMsAzBY5De0+y9nda
Qblk5kh4XQZQ/GHeJ7sTJ1Vj7dV1wNoZdlSQRuENik1w8vZzKV0nOMZ+V+8gnU6ssSAJ5huVpfox
uF3gLMIu80NHmj9N+eF4flvQIEH/kN9qtTqBJHSPw0N7NsT0hG18DrSNktREhppZ5SC/DzHVzSv9
hpj0VRqVi0sQIGEIug1CKVCn94onXH1KigSijO71iql9lh83338+ts3JAHSl0jW7aqzNON9X8jHM
Fvs+Ab0t06Ua1s67oDTWxgilDlNaJ62uUMu8HxRcqrBJUV97FlLIZx5+kM2v8v2uYBh/2hdeKbhj
SfmCW14GC0tLIA1ld3C5pgVVFBGptE54D+ubekCrcneTE+ge6ClRMwtsRzZGtNw0+uUe4gP4jcJb
gDsB4J+8d6nreAfQES4SRzAVkO2xVgo5miqnvJk3axqA/IhcC1iS7ZJKxNiMnpkyvgGrrESWEvW4
tu+YkjMh/di7KfKkAJWOS1XTOpQJV21t7G/lbKq4b8hMZ8Gzl2tdueuRa9qcHJFj/5IXEJllv5VE
byEUTE13QgBcMSEiOZUIQ90l6lI4M7FDJxuyjurxgMLt7kgZoirEB752B45aohC+7Tz6z3OogWn0
mVN+gQEbvHgRqYFBNialfWUkmOiPjeAII4nX/bl8YOwnDcg4UxriQaEEmqmlVBmX/DJttt176n0A
Ao1GuR5fNILIv95griiChKG2793wGAjlApnrItQSt4SbzsgyjIy1GR8HqgWhY+WbpoKXcn4uepXI
8kdZjj6DH05ssix+m3QlcbTvwbOEIeP6Dlfg4XBYFGeCKBxgkQg5CXsqyz1usLJbqK/2DwzEjd1X
OZCiZ1upiBXbqUx2F6pGSNtGL393x7sZnetwHLhanOr1osguXFwmPO6ri+3DgcXMlFkV1EslKjjB
wnUR0HmDdkIwXUROdzhBS+yDd4oy8YVIPRVu2m13L0F/DdFJ7GzzBN9grsbaTUfurfh2R1jzLkyC
ECFx3aDRT24uVgrfcMRqx7u3GSGr7bhzoj4TL+L3rjxB6TILb9x5ge11/YpOVfp7z10PC8vqF+Uw
k8fGlljj/tyZqr5BsMHyiAH8t/FBnjz5KJT26qLhw396PMFARstVhBWsA7PgejeAF1DXHWts/a3K
iRJ/4+FzI+WlEc6+aKxRVlXK9EFLlm/xpw99yWFP6dV2PVkF6EwRJCCACfg+Qr/KRCbVJHVnbPkl
W8vNqj+/3dPpKqLRP8+t3D5CsgRnhs+tUFJJ1nYrBQei6mNXZtIM9AWc2B/SPpqlZvIDRaP3DQ9O
UURAz+sbp5VeZUPRigDpWfnLi+PnVFQumxUTxc3tf9g9vr2ByBqJ6ltwF5dFlzztdBFu2xaL+zpa
Tfg2MaaWHnTlvT+/T7X2+SS7DUbgZ2tjnqfMh+ja1uOrRRqYQc0ZV0hTzLUvY1xUU0MgSer9u0Rr
4bArjf+SN1D0XX9/vSvDAX16PLqv1gEKVJgCAv4R9Uqkmpd5Uff8I/Dz6dAaMZ1lYYBoD2RI9vVK
A3TJtnlVEB80SxnFRE2g0iyAPtaHUBEHksTJhg+7jyGrAH8onZZ9dj5vTa0mXxI9eDTcLO9xhNz/
YLITZM5bZA+te9y4ZGBElWIhxh2ICKCguX2Ez7RoOwZPyQsQGFwjbYEUM0x9grUKQ1uwdbxNw/rW
iIBtxtTRY0gZXPObWZsak0m9jwagCV9q7WZahZ9kd5tnzF5bRtKutAx425nyU0RWsYk3L6QW/Dev
m/dHpX+kWnsQbGSTZvjBQwYfz4zgwvekSps7BuKZqSO6syq0Mhd8dh+1PtAL3/03gLVb/+ddciW3
U68UnLAw4o6lQXlLZPKCKJRrprjnbk1+crj6GfwCQzMfbtdp7xC3Z/hAvthyVbIAyZK1yNcATq4K
yfKvUKOpkGtrant6xHpvFVvmNLDSOYKJUCMS9UJtYD54oj7+tmHzySN6adZFldfqmA4A0q2wv1vn
WECJ/uFT9FdVPlyqeVRQMTQOC6pPsn1oHF9K2XhiQurb0g8fLN8yqZF33LjOA+l84nElWQQ5ldiQ
1lI/L+E05Jiy4EtdnLS0wsmF3+8Sgnb4ZSepMTK9ixgutw6vxmTvITbNA4zjyHalf0dCeCuOuC9M
YLAL4o/3SEGbyMmxEcq4p+EJeIXEqY2z4GFdPmKxw1icWCtJr6Hvidq2yLPvPgxOBy2gVHa/zV8A
m9KcTK8MKklgK+Og8tAOR/fXW36F8XfPtXTlUTwa8cPYQ4INko5NzqyeCHVvhRMZjEXRdiZ5XTjt
PxjbswbT5c9vPhC/R5MriA0FkSegjk9hPumSww+dIGVhSnym6e4N9vcO+yNoLj6POh75iwMhnTil
Vrkh4MUyImDZEYTGCnvtibhZpXrF469KCFI6Qe6BEU5KZBRHWQh4iS2dGQ42HncXpnWm8FWr7Fxj
bvJftls042SP9c5HtiQJvyJ/9FvN9CdKb3znRXHVQPVsmdoIOyHT5XZTNW20FtjlPZI/pHibA9cj
jfvqXPMX7ayrzt9AG14RI5Cr948lLBtxTHcpM2A2NKns3AY4TkWPj4pNAwY5eZU0VG9MlUYRHra+
pNGP2h80LizdAocXxxt0vdLEXCNEquOQyxW0kVaYZlZTFoSmLPn1Ffu9fVrCR1nf58E+PK6ZfggZ
dqPOo7VDHJHNsQj5mXn6XZY0GtjmY3mIrWN1EOPJxxeRfS1UKHmTQUmi3oFbLDVU33O89a6jvq3i
JKxPPxz3IgIW9nbmxwZgggcZAAhJC8PC3EOw8H3vwhMBLZY7cEwBj1XslDYsYL4I67F1a9QqANCm
WOwoVUut9pV58pE+31QtrlqJ+m9WBeIAK0p3HCcsFdkj3rtTvveOQDKCvBvOsSPnQrjTLp3m7GbW
kUdV4xCHE7ef+RkO0HOYT8v9rrM5Yq5cjxIPOYlp+ADZTcTnVObYP6Ll/LO25VHqKVlH/xmTDhpD
Bs+MZiFGVBWDpc5qw1RjvVzINq/DSIFgqUf9q31tsIzr2s1Ru8gyuJY5NU7dLkTsZYjAF1HRvr6a
8Hj8ELShAozZlcuwaaNRb046CKG8UYIAGZuJ6ReSUh10DyVV06m/yNrimrxhhihB2ttIuVGS1UMM
BKWOIV69z9Rc0f4L4J8BYlrWo/qXZbyQYyyciENABmr3mPe8qvWtV7D24lEKjc6vRRJij+RnH3KH
wTAZByrpZMn2Xm5OoILoxyaBnwmqrjMNGpskt/BfmKfHP1mXwizjcRZc4Nl8LAcS9jv+BCL+Jd4Q
I18STojrkFc0ES9SlU5Lf6T1aoMx/E7jMr1epg+435pJvCiPpqiU1p6e4w7yC5vzSAIbqoC1neDk
2rb8BpC0DzeJ7Jz9Kdnw41ePGTxsfwTZ47BTzamcri+Ej18Jhmm6qC4vKNSy6abVvVkGflCa0mBh
lJB/m5ZdIeu27vNfYQX8/yqazi/51RDs3od7VjS2gZi+QRlXZ5sdyiM8BOZ4retIlDlfZ/u3pnJJ
kAA7B1qLZzT+s7IGSQdulJI91XIjUporuczZks5o5Ni+3TTq1PMmacG59RvPkS8r7MitCvZ6uoHn
mD9BZhNoq9Tls19sP0OPUluNGjygsBwgqd6injSwqVMxhQmGT+tfL90BNHrRXmHbo+6Es5TChB0B
i8RYcilkQ2gwwMFg1LpvXcUmFXDA1+nVpScZoJRaR5IptzJ2J/EHdArbfnxxY7yUkyZCiSycwGpq
wUlBiJ+rklY8K+HxzXDA4FWBM0YUSDmVOFSN2AOzeWvO1DtugfzOscVsXeS0kQ5eyj7SBkOwfK+t
tWhAiGBZ3HgZ2iYS8R3V3NrpjijbY+aEva4mxNYxF/7HvbzBAyUoGeb4J3J/gB/KAuyZB3RRPWA4
h2MJYx4GpfCJ8Ri6vF88oKKEVIcE21M2iDlY0z8khKitG/7/KYp+eEr2NbgXMCJqPZsym6qDUJha
x9K21BCd3dYJS2S+p6jljOdiDIVKl36H9cpu++8t91xPo/gMBYL9iOmtVGv2gW8bSjNqGvaZIIr3
dvf3Ht1Hn6ex9eDGgRkOzrsCIOHpZfk1Zlv7I6SNaKAWMnKHDf7HjEHrp6I9Fw1C7BeZ9QFUp2a+
5MJjTAyukZVYy7jQdHmgfJCVkn+cQzp9fjjZm1Ltf1W5A+K6D/zF2r4b6QGcNl96DBO/c5BwciEU
OcG+lUI2wPc36lXDu6lhAQ5IM+NxI25YDsbv6R7CNDmw8sUMA3zv3eFi72YRc4wtiCRed2Sq87Ku
q8IwdohEU1Qh+XOivo3Y4IVLHPMXqHnhdUdLdV6OmcWln2Yr32ZJtLnt7ASC/bWz/5/+JsOPI4hQ
LjAo4zo49f8LJkh04+zl0A81GOeihbxNM2X8/SLZMwKL2e0Z991Qd52/8r6W7kTpFrS/IjoG3boP
M9LrxRV4WdYwqTugiqRSkc1VOnA8Gi+EYVUzY4m6XWxRRFClg+oKpScAKplFxz/fkbCb6aLpmo40
fW7jiJdb2wcm+53I+qBTmt7skXHpbVD8IYupIqw3lNxnbsegWl1f/M2d2qcFv62T8oWqWRDduuUQ
hEMzXGHfo9aN4IJ67tPuZOlPnLuG9xA3US06siwHVvZisXVOvOgNFJfPB77O8jys/RbqrHGT5RNe
iOOFDoNMiRl27TU3HJL5fi3OH5jxWMjWyKyr+v8kma3I4IlkhsVjWUoSfkbjq3at5XNBCls9axKb
lpcGJpBwsanvAGrpcdM9zhzwYbnN1cUKl0FebT9SFp/XUgt6eRbwV7mlZYbPpbFdBJ5s0RSxg7Vy
tlq/HM5QtQNKDKSC/20QmLmUNF6bwoI9N9vgVI7GnGvLb53hG5g/MavHgn56DgbAmdcCg0YgIJIn
8ng5FDsMYGNfatGt0tHM3oaVvenVK/XQkxH41Fm9KALCDafoWtJF6eShfSX0gsDYoUldkqCYkPFb
cKGbxeVGRSqZL/3PMIevxU46bO7bEBw53KhHi06WNcBT4bDSINkG25jhFUePUDdfnthj9pOI7/d1
y6862i42cnkf8DL6tGfLRlfOUtMqBXvhdDMG0R3Oo5BJ7+TkV+l3u99axKad/9lril6hx2iwC22S
cW3RPbbiWoQ4a4qUN5evP3f1NVnqSWnoNdlh7Qp/Rr6mUOBXSKcmL++n2USwMWKLU8INmaPjrpDD
Z8yrpTZMInLBky2u1uazrb0cvMdQKLJ9vcybVQb5quahByyWqEe/b4EB9abQNRhbq380K2tnj0Wc
U4N3NyCrCVimWGWNI4fxRErONtu+kG7yGkWHl+iYcpJxqgCImMJxPqO8no2bMRJFqzgmd9aakWFc
BT1adnmaCI1LS+Xpv7NfS+NOgJrcCzIc1PPHyARQarBN9ELwiRqrR6cVPGjVHdDtXGLmL3AF5u7E
jOBdp3zsCt5NaRy2GdeP22kUUt44h0+h7aC3C66RFjKQ4iGcduK8xE1rw/vS8itiHXJKXjApUQ6s
pGwdOaX+0Q47jSaDrPcb10TuRaVu6soAvGiFlMELFT2CzpdT7hqUksiu1qyyWSJG2d2JavRTG42X
NxqP9XDnhbcNT8fLCZ0c2W/SV2XCNnn5AyUcerJ2V45DaG2D+lliDSrIOqzANC936UzgulM4t5QT
co9gnOENflVpkESFKfeD2+dp+e+o707/6s3uSf4naexXbJ0diNUxZn2Im0nF0M9QBPcrj7qaI2N3
wG6RzUl1sZhLvchyjfqaycP+wmVYxbscZ0/HD/If3OqUpugQaRwVGTxXOyKx3XAGHRR8FW3qjA1+
QFQRz+x+IDmy5cCZo/0c6gbaMhr9RDCbZ/TyiLX/ecn5QDanYsuPNny4gmkFnjJyNUVVDBhntCqS
uAYqVT+LTVvrPhbtba0oT5abDk8V5wOA8ji0uo0k/7uUQK6FHrS0vpZhLg+RM4WSd+RwHZLKKAPQ
TjbAboY3p6RyXovs4FF6NWst2mRny7UwPiOL9yWCp/Ii7RRMiskBGRZCYsVWTuKHaTvLXyB9JELu
YRIqwPCmV1WQmTRNLay20PWyp9A5XE/xTZk3rM5kg/1IzWMjE1yNMDX92zI8b0fEs+F5jzUrYQgx
GbReP/00iVyQ6TWS29r6lnpiKSJrrxNGItLTV60/8me56h/9SLoMTVpazdhXAwsYRnEKkbMM15gM
dWU52OuvZDDN8lyN0aOM95noVDPmmbLGIlnPGRA4Eu4ga/LcDWpV8iac+IDOdF2rdoKoQpy/ct80
m5hTjZsjyBP2dmiR/KWTM38/eE98bTH9i22LH2+1afVN8PAOIGoioegeID0md815KsSvMTM7wdhX
nvJOcacTK3A4FJxZ0c4WbpkxfHF3ESNqh7ALoN7AXKU7hrBxcinIWPflqhqjKT8ZG4/cN4zsgcut
tG6mR7JFHYjUHXI7Z7SetxE4Tgg6ky7b9AN4epUA2isjIZ0rkRhryws7eMxonY4gQn1Z/kN0LbDw
5CxR1PjIIu+OdFmyXQ23Z98aJFTNYX233xejUDwTqZfVAzF/ikp+CArvNwlopbjTbGfQOF/wcDmt
7NCGr2xSoy59DeQyOZREcU51uARedPQBk035GYJSo/ZncHeyL5P5Zahr5uSTRuicq1nOTFaYoa+4
ocTjR7M+JpBIDzQYncbpnDi+5bX4pcUNIyZZ5QA7rsdDdzlNDYU5TYbQEAtg6HmCoaICR6s6iOQl
t6NcPi1BCtbTxzt4p+pdlNHE9CxevWbkVYTxwmOmyT78T5DoOsn845FT73OCdG45kapNTpqdy2e5
amSdZ1zhpnLjgGWd9zt7DECqPAjHnHmWdS1s3yl7hoS7O1SOzmmPFjkTA4mpI5vJf63f4EInNXAy
OYpAUy+lNxdrFEZFq0DB3sYga60miKWR2yhPhLTT1HCVcxq8DiVCT3T5LQewxk/0QwWQizEqH0L2
Tokcf+i1LZdDl7GeBZzM13uQUjWZVItpTlbj/NTyxWtdDtgnkjD97w4Nhm3rWsGB2jjU3C5630km
cBA15aiaqEqMyuK3/RH+Y+m2WzF1esb2IlkZJTVcnxHIYDYs3XXYB6oBacgaPbIoWccjpFM6uXt/
4l//+D9Lhf/u+4EdlnHHM87HMMBQI453VpSmJ1/Uq8OIG4Mq1jY0elFrU6FGlrRGc1n81IZJkiHH
FpW5ZdgWSBZkWkqwCZ2f77+z4tbHvfVRswK2NF/3E+GiBJxmtaAxOBzw6VUd//JgFx3Iaq8cMa3L
IBfer/AHyFBT9+CQe2BKOOG5daHh6OFql5IwFV6u6SkSrmIMA9cdtvqSK22kS44RRBTBazhcbgkh
/J3Sk1PAGjKwwtZDqvMIH2963Z4Hi5MZs5iw13lGJMYo06mnfyS2KwwSmLLIb2T918ltoqQur06s
xDJojbyQPUrU8YVeINj21S6V2Nw5mDja0CnhIosxBKrCp970gfs1aoUA3/O1uFLlLdU1cW9n7ih/
bX4i6wsnV4OOc0gy51bYdl6w5c2xaMAryR6GeLsGA463LsJP3xNZxTnnAuNZ98SmTPt689nN5KxC
MricnDCjiXaVMAlhtSftgN3ywpf9mDW4dhjqHVvFaeyTpSNpFSl1BhB53VCR9TATaa1aOMI0z9Po
ZxKBZ7FRsyShGfNgFB5qauWMQlpL0qivNObv15GcO3tzQNcKJJZYGook/K8l1UA4+mL+lt/UmRLG
djq5//2zK77vBaTTTNS+LbyF6baiP+1TRQsrST2Z4kiaN8U1Axr2/CVIugxFWTMaAnPxlTC19qyk
KHxxTNpMbgddepUrSu2aOOlpyo0GKCKSy/yoIB/P9/48r5I1QqSANUtQ1ajfFJxeWJ/b/P/Z63cd
UI/Dub/3BpXllA1nd5vlCPKnmIJMIC7hdoEdXHqCN5MMy45HJd9R3Cg3DErPkq7FrLal5QjMuQoa
J1MmU28GQ5b6NjQs27cqWFwSwg/JZuI2862zneOQzun2FxRG5K1rZODYh1AcQ8C/jltHV2cVYIHS
OETj68D5eXDal5+PdCfyF26Q6pNGUExZW0E2uT1bT6a9UTAUcRhnwZ1nye9MS02Wh6SiyYddU7Sa
IhLXTd5d532BGQgt1mXY/8HKDXmQhdwJROq1/1a+G2GNB0nr89x1MfjyS8lvDk792tQIABcuRjBA
slZXE3y2b32CDIwnixZ7X1sR2GDvZtfbdx/FqNpNpuSGbevqIbo/NiCjlRxqwVLGmuwILVWyxOXC
3wXgDPfeZDrw045nOzMyRNo/6dwZkoxkY5WFkf4r7Pe+3PlMf+4opndY0FtohZWHJhYMHqFYVL3z
7Shs5IXG68gHkaZ2qA953WD0wV7q8KFH9P/4LwPr+C4P+4RR3dLGgSpkcExkwJSpdB3pMGmeBE2o
+TyURqNtaDeimL19UJMM90jC37D3i6L+CYQWlUhrVsJxV0aLc/WCQqiSwLq9kwhjvzC8qkqK+ySU
gjGXhJ6PmDnqidMAVeXwDV9cV+EcD8WR4pwoVZcgiorHwGpaHX292GQ59GrgJGhhy9fB04It0fSz
9qbIXbq3UGN0Z3v/VSIF0cfaj3AHpl/CXYgjmTQAQzRAD84tWQA8Ng3eDA8BL1GUCOCRzblT3dG9
+ovIjl5roW/rtf9sjZMKGl13JFbJ8Hf4HAFlWcR394lWNy/ZUpR/wDtLV6bGEJuaxV6/i1eNSKFr
CeSq13doa2rZ5wxSfS+hZo87d/9+Hf0V0ML3Vr343Y7FDuaAo3+qgkr6KuWtFlXuqEliQ+MQ7yG9
/RcK9JOp3WJTUe1F7oJo2ZYigQ2Zl6VihbIOVt3+sL88D9KP/ARKv9CgSYhWc/pjp9yJJ+L/YpfO
U6D9soXjq7lBFD7uyCIU4JbDDa0kdQr+DZ564t2FYdcwugg4otIrJsxagYkH3MIs3rpd3N3vvxzq
zqtaMl37U3+Y7zroU+dTpscM5FzqUf7mfl285OjUPBs5V47j/3+dHzozqAW4ZqIqjOlPNVmo6Qls
79IXRfB5c8QuVOl+NOwzF+UOjg3t1lTpRLrUdbNe7xTgMGhH/XA5f0mUBXKeQ0vKS5c5CfHlet//
kiKB9gbC75pW8Y3YmXA/7/M9/4bQ557BhOM2cV34a9azcBETqYjCYDl9gs3+8zGS9gNT69J/NuMc
hfuVkarfRWpqqiQG/qPMCWyg0PGn5eEXAA+1rBF6AUSrWseKtgRM5gQJeoRhOSKh0an8rcQveSr/
FWXijL4TS1GjOmD2Of7xLtI/m5M77WqIVV+P5AVLwFf7LMMFNczrn6Sk8numzTEPTYwwYHpbvExm
cIMhpCbCK2/YMQ6rVFHtv50Shjg57CI+yZxkMirI6c2jo8uADiux1v0jFZyGa+sgUt44idLgN0zk
Buv2RypGBn0bYFSS72FFnz4AU70dLFxf01WA+t3+G1wuIBNeDJcr1+Nr7F1kxhogeA0xQ7E7DDQn
SbFmJIQmn4/hu9dpmA4VRXXcLSPNy3Mlmog8sLV5v9oerFCDUqb3Zc+Q9Nk4wVK4hLLt/BY22gNJ
Y5a8SE8o9CDwF4mFL7vVMALJLYEQe8U61wbmq4smuCn6tVg86KL0b03fWZnjgAGjhRNpoiyxLi27
xGKbO7EBFJKMo4pOHFU3E7dzrvOoNtACEhuymOP1/xMDaYrGoagHEdpdlPEaDlaoDIwqIWZQeOdX
mYaIiti7jAFf6cT3bom4YWlrZzWmp13CuBikyVpUhdvF4XojmLIGL45Qcc9tU6IVTtr8mEYkmljh
tzAkdb1Kn96E7fnitIDhP3PaRjxc/3JoulKcpR/WzeObLtdIDrwtOzG9PNVaE6mCstzt83jum012
IKXJ+E1JZrXMKOV/epvIbwAZSaksl1tTIGlA790aDsCtAoWrNwCIFgBUxCbxxISz4W0SX10/ibUf
Cg8M4f/jWcP0TNC+J9qT5J3ORqd042Ti9cezKR22FekCPHDegFKrmAzNAcQk03HoYxZcr/zDrERV
CuZemlg5v0fVGs1VWg2gta1X/T827Vs+yLviSFDX5HhkqgsQKeL1Bq2hIqzBHqgACoWipIrONOyh
HDk1lcK/opCMKedENnX4BgXtZCttfeZ/NiJh5aFNEi38kU18rQjv6OpJdQxDJdWuo116Trh7wwzn
HvsSrbwR/qI8BtitkuDpsJxTBVapmheNN4qtWoxqsejr2d2vcb586vEY+RN/ERXzGbZwGks8tKSA
4c+oe7HlAFFVejIiaIL30m3qyf3d6zfqVSsqc6QtV7tvbAlzDUJh+SRRTuGyFYVBLejIt0Y9EAiO
5t17sYRe4PtRqqGmwluI0lXrDleY2YVAiDn+llkzT7Y/pBDh3ApJ1NWOQyjPS96Z7cFOIVvF86Fw
7kaksPZrTfamnrIolZzb+Gk6P8VZ9yowIUdomw6k5pcTXvOoLHeqrwfkB3nPdEYdczJqo1mfYLN/
w1Lk333t0M7GF2SfXGXJPWmHh9ylO7C7FpawvH6Swul/WHjE+l0mZD1mPRWoB3LoYFNQF73ON+vP
cM7hdmDB9Xw2HYSNy8EfO5niU+eL6kYVHuGxCS00ZauerZPYsWR1+dRSqJdXHjM2kddhxbFGQ5VP
X/UomxH8LNIIQHuOraCJ7QyKWfLLgpfpgNFW4FsIKIIg4WeqsQETZyh3AL/7xuxYn89fQk0Opu3D
HKMEojstT1dcq3O29uUU2f+NpawT04NphydmuFiMftdTUYrVHP0slCHLOsug54rvzLUNUhJ2oZPW
8gfMeCgQALdDXXtjLNZ7DxqREMjoscrqalg+EjsUWAHgx8r5x3BVwvBJfeFc1waxGto6kR2ljCvT
49nCtQd482gH9dFFQ5oFvPRmIOqSFqJm3xz52Q2qPlig7fX/P5+YvE0HzATXJFFgLHjYovck/E88
pV+kqDze5Iw1v4sJkPDsdiOnLS2eSBd+x2bWs7D4afY9TZe/5y1hPg+ZX3vOYbFBfFazKWqYknfH
NA9/suEqLxMSs+xKA5kNbtH/SZ3+zBr1wSURVekDxbUNj2DfJqQqkqGhLmqT/yISALt2aCh/seZG
6bsATsYXAbx868RcknEu/34F2Q7TmRlw+dEqLswQuoi85IdVsLdAEZmHxe8be1rgWkVoIh+YWiVp
bp8W8ItgABCPrAPyG7jTVX0uULq6fEEQh9Q1hxFn25n2I2yKzj4mcqz9g1HqtmssjtbeaAjJrRKK
mFxhNurn0oHXgwJafXUeUNSd3btkzRe+jhLVaYmOYVJH5weoKRdldSyPtFDOm8bRAgFhhiSQ72FI
uqVkky4dEIpK76se+d8VFrjFs47CHCt5OF8sCzMVzvGH3hMrSWZaayteXtWPtTtkwxjADAcQ0ItU
qqJsarEFGwZziZQKfM6pT4FILZCRn0SixHOd5XwP2GnKPAvCUgo0UYsINf11w/7bkEsJvtBlPuaf
KXHfSGvsFaklHxZ7doUpL4y6anX3SiOTDlk7bqK9SDQM4z8oxt7avQ1/dwAERVacjAkdUpXTJwCM
uCRXsG7FC6pjsymJ0EmWB3ZmN+L4A37FPhTcbUbMVd4XAZDrF9gUVKCSSnLriD2ery226jlPnKmu
qyIkhklXBgNSSiUUzn9vbB1Dnwd5Q5u2pz80+WLZdTahi7+zLPfGU7EI93fvzrS4Sng2B0HB4D/i
W8ezdE9lEocWN2uVnS5wqXP1z+Tmn8c/umnFo1dD0tqFEKnkN9wEKWM0uJMz1QY93UvlFoRy0mi9
GpKbNMlrEBbFxmk/EN5sxhcaQYHgX2grs4fEMmP/eneLygYCtG/5W4nUb5fqJYkAJq9bnQpdwbTB
4yQG3tH3oJFgl5RfRBZh0ZgzhBy+hU/1fYCSuLJPJ6JjOs+9wODygR7N8rraLnL/aRcsjuL+liHr
A0J5LkKfzCeysIE6WRPr45ExoQhRq0491KdLdfCyAluf7oe8tiBx1EhHZiCl8Wit+8Iy3GcTY018
gzZ0zDwRMGFy8GXNUzCw8WE+Cd3+D+//L6L9jyJPSLI9l5Vuy8ZSMvzXVKqtgaberL4aDXRp8V+T
V/s07vPpjxJ760qMXLQAhawJ2TZoBq13dz/OrBouPcKOY3bTEQqBoMldzV6YTCHdKbG7WwHTRF/p
G2SaDt2qkSS3S5bJ8WMUxKhUav4a0BvwHpKjCuoyFDVJOFUsxVqogDaCVKnFDf9G7dmDyitvF4Mk
2mOBb5W4zD8XUggj0upikY9qPOnQyH4S46UDnxedNnHO0ZGjV1K4WypZ/dpAQZF/KN5IjI1/3oM+
UEihOKFIwIcwSY7l0ilyMKDKutXB37ZaYSqmLIr/KCV0ZjVX4S3gH5sXeC7HZOONFVLaioPramIf
449MF8ZyBO//8Qlgc6Mu8C1zn+i49jhKVJBdWC+f79273FxDJ5BFxB9l5Sj3aOrUEAS+UK19yOCm
gKDgG2J1dWo++kiCyeP+KUbE21DjSc6o0uhbVs31ehshkENuRc8LNKQSxI7VgJdTZaGCl869ghZH
MJjHOEa3Tvy+0xoQHBrSwc0Z9crf8D2F4tJ+bcNj2Zpqk37XkUeHyFWPYYuJ+/lQZzmRjPe2A6VT
KgYnHQQwJnI96m8OzoXto7CArTiQHJyHGvwt+UXpq/J7zud9vbN60RgsXK3aAS/Gh72ytLgaKdsB
GZYltgdj8BUhib4KAuN+A2tmG8Tgquv+5TpsFJbtTYP/d+4yeUyinXEGbJ1vbNDYSIzdiWB5WlnW
OCth+QEpXNACPsPv0ijM06Jq4RjFmQYS4I4Ek1slFR2F6kARnxVE7L+V+QQEg+qP3dcLWUBr6CN6
Es6o5FN7WY0p6NRV8JYzD4LJOVBtxJV7ptrWG4LdT5Kk6fBxiotkHIXRW1HczQTmyKWsPQ4CUTOq
WPy7gshHzfY6nXLzSnim3+0xrvAWAFtKhmPF4GwAWCgpU1LRyu+sTt6JBWWpjHHmCJxXsm2hCl3+
hvNJTrWYPuCi1KeJubjTJGVHc+FfoJP80gBr5FoNMyAV29DlqMh1J9Sdk72kFjCfuI/LdFk1KcBo
W2iwNWKGV3JdMIARrO0mWDdM9rWNhQfZ0oCh9+nu7YnjNhsVrG7ZVr/9cjcqPbX5uSm2f1Lpvrhu
zvVwXzJRkbqC4WbrZP5j+FsXR7dWQeP4t/YwzXxI6FBlsrWU6envNp9KTuKCgRWglWA5phKpIpMj
UP7EtLKShNWi6r768rdJIRXodgtFlW4ezu/gZ6vs18stOA9omgISZsUkpqmAoe+IALxmFMzFQ09+
auQFwT0nRL1rUgEU7FT46pmJCdcHshlNnCiLbjjsieNbzuvyO/EG4W9CyDdYeBMN2ZhN1zbQ4L0k
2Tv+2gGjsliBTz3Nc/dC0RdiEEth6rN3sTMqUk81Hr+OVhemGqvA1A0e/PDTw+QyKeoGthDtHsLM
49rCk8wtlMN02ElnoHYGKXALs3OuP68bEgpRZyNW0/o77pRnDgzT6X4Nt0rrT3yW2BtwET1jPdap
LaiZFHVb/u8wKhQDMrunE5+kZNkgPScWh+F+B+QMMbd5gdkqDRSz5MXUgKWV1M4vfuRTraBYlMCJ
HmjTsCIPwwITS4V+eHEfvg4r59PY/xasHAJhtbsoPprEjKx/WHH3E9eNklO/YkZDe02B+7OETZrL
tgCAP24F0MOUZGaidA5Xlnwj9rYH2+IzSvJ2REDk+wBjcvlPG4H3bdUkngOw1yW3pO+luIyLxQSP
A4ngcSB8A5WdqHIrWPK41mV5E480AVGRNhMTLd9oTquQ/155ITZk7vo8tRLMYk3NCzAhxI49wySJ
IR7KfC1+1iJupe1qVoe4mzwwFLCcDhe/iAix1jqRsEobgIlG0EOP4tJJhKB61du8pgGkY0A0NvAW
K7XRpUB+qRahaOpSZxFaucRGM9N65qU1aJ9BPdiZv4tVOugn2+uSKFd3TFvmo2SLBOf2hhwxwl59
6GLd8cfOx7JPJOZpx0xTk0eylhVqWYq+9t+RzpD+sSbQCLAiYe0zlfE+wVHnqp/rsHEG6Iz8zCcf
vFJ3VmVKXuHcu8FTHBMaIedDQ1aFIznQkdS+WotovYO6FfjBYob7YCnMQkGMqHFeq/RrKWBE7fxi
j0aXYlqD8O70Kco91retJgVdv9CdIHBK8X/mge3d4JWAeB49Virj5y0XrfoXFn8mRfviziy/K14X
U4jHCXOzqIBHSgmODCloILv3SlpLoCMwykJ0OoYKMq/fGKmAq6hvbkMjKxqUzeAOcnv5dYYTW84l
9XTy+yF8B33Gtq/eH9CDV0EdUnDSOJSWHNSY9oc9j48jp5bTKWMcEm16/lx3kkdjJxEaRkiwpRXi
iM5tNc+6UqWHGgoUxJ7ksUZYWyaBatKdAcWV8o0Rt4HGTPZjFp0COgumiVC5b/n6w9YSc4HEqCup
9jVATnsHSAWjuOlxmK1IgrW6rhsXiY4izF5ga0PQbW1/aZ0oVOmOajGUEyV8Zt2zkCXZKIJZdhtE
L5jMcEFekNiSm7uyMeskBVs09auHafS+rAaZLeBag1R030nNnSEzMQPHbmIlZBkfoCAkkpDAA8d6
irktj8oHvWMY9A2RTE5iSqBNuLUXc7yzI2UwEnDgWYyJ07NAMmRBWr5fOJQrRSZkkNnwQMBY6ekG
MYIPOK60/ycZ3+7N/PWycn1scC2JsCP9Dvc1ZCwJ8gjiOsw81K4WBo6V1NF7Fq+r74wRQ6sGbMwr
jGaJt12ORhl0UDHQ0zHhTjWztB3BjVvtMmcR96aBJkc5OLTUmvmqNmposkavdDBMH7PrI5CuoZ4S
lLVwKY4Y2CsAht4tj8CZ+ElbljOC/So8Kdkih+VH7Vc70D6UH8eK2AdNVhVVCEA/yIJjX0KPy8/+
EyNGS5MhMYKaEnJLFHq96K2V+UPBQI6pNqB5cw8Z6bdNagd0+oDUxu+6s6TXCcj787PLUKKwQzWm
k4mp5e834O7CMGD2/H2NoAvZWsTizOm74fpAk2/B0UNyjOLt0r1inLa27CR7scRdbfQMpmdZ7nmr
Wuu+6JcMBf7Q/B2SSNuOGlCIiwBBC5x+cRwUcz26lZqJ+EtX7KNIUO5GwgZZe6enzVy/9J/POokM
RhLsKAKdcw8HyFL5TXOK/gpb/yUsnbDJIWWL2WLieY99SW7DPD2sdgrn1l8uM1RauoKuXPOXR0qx
4I8dObj4/M59v8db6xvopv9mowFDxVgqG6gxo+PCERlfj5mAdNIOEJLszGgxHwuZ8HetPIAyQH1D
x7R9Xtye2MmqWQlCbaU4RzsrG73hEw0Md7y49Daqgm7hnaSbFfY/ZMQLqzS+N43vQFspZ9oGfMXb
FUITNqQcDLSwp8cMcrwbFuXnW4lqpRmqsPejQYfQPpBqq/PBfMWpmZLOEIyOiZt4QqlnUeTz+em4
/vmvhvXd+TAPRBrMSF8v+kLeIJvgip1Mz1Qstq8M7MshXH7V9R9g8qs4ksWfl26EgT8grYQ/5rYL
zWZ3f5Quwc/HxGaysjUaSoKB4VhNJv2GBUny6fDAarLHHsHplHUj/DjBv0HT3Vx38j2K/Gx/H85c
aiB+I4DSpPtJl/bR7K+Wq31B1sSvuZTD4OzxWRlcOVXz9b8af3qaOwlBYisHNM90mLWjNcEn3Op3
gTGUv+MTFtakKaLDYhOSLr1MsqsCm0Lt8H/SLslYubipCI+I+dhihPvyyqJDV1GKhxK16fG/RySC
nodo2VkkGBcN//gmWFg9vTlnTq0JckmulssyVMv+h6Nuh7HABdw1CQlkLjq8uonIV7oEmNK2laY3
Olpsa52yw0P6gwXTQ3jW17bmHKSLJ/85sjo7AiT7/2uZ/whIxqyDryqzlyU0PWb7/TJ2fJmcYEq+
4u91wX5DIaMmVBqmQplM9YV7Q2oOo0ibQksK/VAKjrdLNIXEtcIWp0tsOduGsFE9svJApLPHwkRl
o7W+tyW8X3PkV6zeFdH3KO+a0O8ZuClBH2MebuJyQtPiXTi+a8x/iBPiUbKjHx0qox1dQYiFwtVw
z9affgGag4bTsL/MOmsttI7Fwz1izekPI+RRmRsVmmuW2FMRlAbF0+0198zJh8XryrrSQEKoWXES
24L5Aw6TQZxMjpUP0cUmUuF31C/nmuC2ExTgBOhB4heRJoebPMf76GRtMhTDYHK62vMmSnx21GQQ
KE6jjexjEJCD/GZEkvpEjh5R2UyNS0ii8QQ9/dAuWT0kPS90sRuY4K9LTykc96gH/btzNMlaDFR7
fjTlWHPRfkYu4H4R60MH77XbcuzoQN/LzIcBbT7/w69p8Ae8/miPmmr/0q1moCBEepMuJCQIVEfH
OFCSLFL61PIqwFdUZEwNwbecHpzkDbMtqHnOMReY1sC4Kg6Tj7+iJCxlLkf0tOUjhq3sV0WVokfA
X/l9IbTGNKuTuW+vJmnKAHS+2KqRKuz24pJJGsleRBQF5uYWY0/zRBi5HG3duW/0dKotB9Ou+wD5
2uN6S7xQxowFB9myJBF0bXSLe3IEHTEBByvNO5eMJ+xhWCZkjCCQ79QP+SIAyv+l4HP+ezc3cYih
d+buTfI+KxzyEA9TQ2vYB8qG3e46kebQCcubVIzm7X5MmObQjpa0ZJGUW0nHlbWWNdfayKrBbK5M
IHTZLB8JeGXLZ7GuFL11Vy3JyQ4ici9db3D1qVEQiqX6OhbAOFhHyHFs9CCWXC+oNmnDGLjqlMhs
gtW+sMAWnXqNZ/3ZMyYWS2NmMAR8Ei3nE4mrB96zYnG4XEgaHai69D8dnMsdYsWGQjLh0xxJm9Wt
Om72WApqW6fHbv60izedw3ihL2EAnweBaPHyt3JzaZ0/dnctiI5+WEbY7GmMi6o9cCs61YwfoPLl
/UaXtJKTSDv1bQSPYaiARypochBYKOOnS85AC1VyzVkChYnfuHHLxl0qf+DWb6HHQpc4L3oHYy0I
JpkMOMK6cz3dCpIvLSnnuyxmL4rsiQtyKVL5HZIPiVAfO1/cEmqcFLG4LeH3hdAK7PbucSbyv0GK
87piBIc+nn6gGUKMxvcfAs159K+Cow0ZOrhdnDqYHc/s9o4vBe+iSnrDRMdj4KMpusz1xBbJbPwy
bBXLvnHibXDP6Wvp4DzqBwvRNJjR0VACghZjVNuhOT/Yv4VI4xfN9kufVgrqkaxuFsK8DDCi6ZS2
TVIv+TP/6Bi23KWrnmfCRMUW2S7pVDWtQst7ppFKHustaYreD7V9RiTKXyjUWMmfuby2ZQhBKRvI
l8YI3dskTGNEM9FZc0e9bN1Q8R6FYwFYxb7D6qCWUpeEhxh3V8eCJbmA7T8epDApFffMbD66GebA
QbFwsEiMt/oP+2GH57ehFt1z94o3cWJ3PpYImriFZBmBjCfJW5OlTZUVOPEhsn/zfKbWpCxKFoIv
6KndiVc4vCnjyYfwWPngA+rsWG1KRednXUPcAkFqTMZDy9dKdm6JH1dpwm0k8cHCWz1i6F6bxFU9
gqqh3z8mRHJAPugXK4k/5/JQTdLmzcTqamJ28mY+ibBxxWt+CjH4t/1BHFJlZna9PG0q3mA62C+g
k4VOUDwK6K57Uyx7j9xFhZPKFKhleE/QN3fUK5bVtba2nPryz8IRIg3ywUZcGdWfB1g216i2+mGm
PVpGlVC/t5aPhgWtE4jjVagKCaB4iShIjBszmhpl9hQ5uexKMzpycmHp9pX/sJ7ZVyreZyWmQ23L
fq1lnrR9UecNSKR7MNtYomL+1NmaPHGyE0f5mQ7dhH4sYZ57SJB63Rs0Vhh3lmY4ycS0T17Q4WHN
riY/7axAHzP//4RJ454EZXT1UsrRRIB763I338pjy7pWWr1meO8IeXtCLFbAoQd6OkBxRDXsWQ28
gQ0GjNf2Knq4etnWcdi9SpnQ8mDlHFjEfK5mY5Yzd9tj3M/qwtK0h3NM4RTxa8j+5/Mslcv9terW
JjmIgoTIAhEdsiabsd7e2qGfwaEb4kF9iFcNZ/WL97MXnZ4e0QmNzPgaU4LsmI9/R2TxMHCZD8Hr
rxz3cPfN39EKKf+0w7lFG3X9JpIGJF51P04TNJVowHlzFy1JKojQB6a8Rt4uD1V+F9Q0hHim9ogj
tAXMpcFMZMgbUOUjXFag4ApT91kE0kd6VV8GopVfW2KBuBf0MA3VvN0culvPKoE+JH+NWx93qwog
I4eBzBrs1Rh4WoR61Q4a26jIQN3DqHTZnWYZZjD/5Cqzcy8KksjzZUxjwZ+8mQduEFYn3BUdeIax
0FNzYDgVI524U2h7I6Iho0BcLhB8iPPov9ymz0IQSUQfS5z6JxYKoTyCFy/FYRkC7upkgI1t5AoJ
OFNGSKku5p8GM66Z3a8oUFX+Q6j87jB2wMH4kT11L+v62e5UxAmYivxY1Wc2HPfrIBFkKuQ/p8NJ
PQEXKElTvl7MiwCZIgu4fQemQ3zsw+PUJedBtT5f+ksV8BAwJN8VMtXbtkY927hEVDkSxPq0FIFC
3ll+iIES9a9uEwA/bHX6mVIQQH64Zs/10BD5EB+6DnqLh4bxSeEKSTaC7uho61yNepyZ3qF9TLJU
AEfthPmrQM6d7ESD+otqnMhnEMgb1ZFw627H+9EmXXTB9fsrE1Dv1PE0NPaAOa1a1M4jDbUN52/K
pReJRPaOT65QPn/zLESpjw3lThSM1xV55wX2bKQjP0WnW7hY0v+yqLzTlvLb0gquyw+ZsshMwr53
rRcC4Pgny0nzNr7KeWrFY7ln6lgVkBNvhPvTkthV/OkPV2PMurjvGl+Ug6aRnd2YmpGIaUFBfZWh
n1zJBYUL9alSMCcv+rs=
`protect end_protected
